module emif_ddr4_ddr4b_altera_emif_arch_nf_170_3eabgiq #(
   parameter PROTOCOL_ENUM                                      = "",
   parameter PHY_TARGET_IS_ES                                   = 0,
   parameter PHY_TARGET_IS_ES2                                  = 0,
   parameter PHY_TARGET_IS_PRODUCTION                           = 0,
   parameter PHY_CONFIG_ENUM                                    = "",
   parameter PHY_PING_PONG_EN                                   = 0,
   parameter PHY_CORE_CLKS_SHARING_ENUM                         = "",
   parameter PHY_CALIBRATED_OCT                                 = 0,
   parameter PHY_AC_CALIBRATED_OCT                              = 0,
   parameter PHY_CK_CALIBRATED_OCT                              = 0,
   parameter PHY_DATA_CALIBRATED_OCT                            = 0,
   parameter PHY_HPS_ENABLE_EARLY_RELEASE                       = 0,
   parameter PLL_NUM_OF_EXTRA_CLKS                              = 0,
   parameter MEM_FORMAT_ENUM                                    = "",
   parameter MEM_BURST_LENGTH                                   = 0,
   parameter MEM_DATA_MASK_EN                                   = 0,
   parameter MEM_TTL_DATA_WIDTH                                 = 0,
   parameter MEM_TTL_NUM_OF_READ_GROUPS                         = 0,
   parameter MEM_TTL_NUM_OF_WRITE_GROUPS                        = 0,
   parameter DIAG_SIM_REGTEST_MODE                              = 0,
   parameter DIAG_SYNTH_FOR_SIM                                 = 0,
   parameter DIAG_VERBOSE_IOAUX                                 = 0,
   parameter DIAG_ECLIPSE_DEBUG                                 = 0,
   parameter DIAG_EXPORT_VJI                                    = 0,
   parameter DIAG_INTERFACE_ID                                  = 0,
   parameter DIAG_FAST_SIM                                      = 0,
   parameter DIAG_USE_ABSTRACT_PHY                              = 0,
   parameter SILICON_REV                                        = "",
   parameter IS_HPS                                             = 0,
   parameter IS_VID                                             = 0,
   parameter USER_CLK_RATIO                                     = 0,
   parameter C2P_P2C_CLK_RATIO                                  = 0,
   parameter PHY_HMC_CLK_RATIO                                  = 0,
   parameter DIAG_ABSTRACT_PHY_WLAT                             = 0,
   parameter DIAG_ABSTRACT_PHY_RLAT                             = 0,
   parameter DIAG_CPA_OUT_1_EN                                  = 0,
   parameter DIAG_USE_CPA_LOCK                                  = 0,
   parameter DQS_BUS_MODE_ENUM                                  = "",
   parameter AC_PIN_MAP_SCHEME                                  = "",
   parameter NUM_OF_HMC_PORTS                                   = 0,
   parameter HMC_AVL_PROTOCOL_ENUM                              = "",
   parameter HMC_CTRL_DIMM_TYPE                                 = "",
   parameter REGISTER_AFI                                       = 0,
   parameter SEQ_SYNTH_CPU_CLK_DIVIDE                           = 0,
   parameter SEQ_SYNTH_CAL_CLK_DIVIDE                           = 0,
   parameter SEQ_SIM_CPU_CLK_DIVIDE                             = 0,
   parameter SEQ_SIM_CAL_CLK_DIVIDE                             = 0,
   parameter SEQ_SYNTH_OSC_FREQ_MHZ                             = 0,
   parameter SEQ_SIM_OSC_FREQ_MHZ                               = 0,
   parameter NUM_OF_RTL_TILES                                   = 0,
   parameter PRI_RDATA_TILE_INDEX                               = 0,
   parameter PRI_RDATA_LANE_INDEX                               = 0,
   parameter PRI_WDATA_TILE_INDEX                               = 0,
   parameter PRI_WDATA_LANE_INDEX                               = 0,
   parameter PRI_AC_TILE_INDEX                                  = 0,
   parameter SEC_RDATA_TILE_INDEX                               = 0,
   parameter SEC_RDATA_LANE_INDEX                               = 0,
   parameter SEC_WDATA_TILE_INDEX                               = 0,
   parameter SEC_WDATA_LANE_INDEX                               = 0,
   parameter SEC_AC_TILE_INDEX                                  = 0,
   parameter LANES_USAGE_0                                      = 0,
   parameter LANES_USAGE_1                                      = 0,
   parameter LANES_USAGE_2                                      = 0,
   parameter LANES_USAGE_3                                      = 0,
   parameter LANES_USAGE_AUTOGEN_WCNT                           = 0,
   parameter PINS_USAGE_0                                       = 0,
   parameter PINS_USAGE_1                                       = 0,
   parameter PINS_USAGE_2                                       = 0,
   parameter PINS_USAGE_3                                       = 0,
   parameter PINS_USAGE_4                                       = 0,
   parameter PINS_USAGE_5                                       = 0,
   parameter PINS_USAGE_6                                       = 0,
   parameter PINS_USAGE_7                                       = 0,
   parameter PINS_USAGE_8                                       = 0,
   parameter PINS_USAGE_9                                       = 0,
   parameter PINS_USAGE_10                                      = 0,
   parameter PINS_USAGE_11                                      = 0,
   parameter PINS_USAGE_12                                      = 0,
   parameter PINS_USAGE_AUTOGEN_WCNT                            = 0,
   parameter PINS_RATE_0                                        = 0,
   parameter PINS_RATE_1                                        = 0,
   parameter PINS_RATE_2                                        = 0,
   parameter PINS_RATE_3                                        = 0,
   parameter PINS_RATE_4                                        = 0,
   parameter PINS_RATE_5                                        = 0,
   parameter PINS_RATE_6                                        = 0,
   parameter PINS_RATE_7                                        = 0,
   parameter PINS_RATE_8                                        = 0,
   parameter PINS_RATE_9                                        = 0,
   parameter PINS_RATE_10                                       = 0,
   parameter PINS_RATE_11                                       = 0,
   parameter PINS_RATE_12                                       = 0,
   parameter PINS_RATE_AUTOGEN_WCNT                             = 0,
   parameter PINS_WDB_0                                         = 0,
   parameter PINS_WDB_1                                         = 0,
   parameter PINS_WDB_2                                         = 0,
   parameter PINS_WDB_3                                         = 0,
   parameter PINS_WDB_4                                         = 0,
   parameter PINS_WDB_5                                         = 0,
   parameter PINS_WDB_6                                         = 0,
   parameter PINS_WDB_7                                         = 0,
   parameter PINS_WDB_8                                         = 0,
   parameter PINS_WDB_9                                         = 0,
   parameter PINS_WDB_10                                        = 0,
   parameter PINS_WDB_11                                        = 0,
   parameter PINS_WDB_12                                        = 0,
   parameter PINS_WDB_13                                        = 0,
   parameter PINS_WDB_14                                        = 0,
   parameter PINS_WDB_15                                        = 0,
   parameter PINS_WDB_16                                        = 0,
   parameter PINS_WDB_17                                        = 0,
   parameter PINS_WDB_18                                        = 0,
   parameter PINS_WDB_19                                        = 0,
   parameter PINS_WDB_20                                        = 0,
   parameter PINS_WDB_21                                        = 0,
   parameter PINS_WDB_22                                        = 0,
   parameter PINS_WDB_23                                        = 0,
   parameter PINS_WDB_24                                        = 0,
   parameter PINS_WDB_25                                        = 0,
   parameter PINS_WDB_26                                        = 0,
   parameter PINS_WDB_27                                        = 0,
   parameter PINS_WDB_28                                        = 0,
   parameter PINS_WDB_29                                        = 0,
   parameter PINS_WDB_30                                        = 0,
   parameter PINS_WDB_31                                        = 0,
   parameter PINS_WDB_32                                        = 0,
   parameter PINS_WDB_33                                        = 0,
   parameter PINS_WDB_34                                        = 0,
   parameter PINS_WDB_35                                        = 0,
   parameter PINS_WDB_36                                        = 0,
   parameter PINS_WDB_37                                        = 0,
   parameter PINS_WDB_38                                        = 0,
   parameter PINS_WDB_AUTOGEN_WCNT                              = 0,
   parameter PINS_DATA_IN_MODE_0                                = 0,
   parameter PINS_DATA_IN_MODE_1                                = 0,
   parameter PINS_DATA_IN_MODE_2                                = 0,
   parameter PINS_DATA_IN_MODE_3                                = 0,
   parameter PINS_DATA_IN_MODE_4                                = 0,
   parameter PINS_DATA_IN_MODE_5                                = 0,
   parameter PINS_DATA_IN_MODE_6                                = 0,
   parameter PINS_DATA_IN_MODE_7                                = 0,
   parameter PINS_DATA_IN_MODE_8                                = 0,
   parameter PINS_DATA_IN_MODE_9                                = 0,
   parameter PINS_DATA_IN_MODE_10                               = 0,
   parameter PINS_DATA_IN_MODE_11                               = 0,
   parameter PINS_DATA_IN_MODE_12                               = 0,
   parameter PINS_DATA_IN_MODE_13                               = 0,
   parameter PINS_DATA_IN_MODE_14                               = 0,
   parameter PINS_DATA_IN_MODE_15                               = 0,
   parameter PINS_DATA_IN_MODE_16                               = 0,
   parameter PINS_DATA_IN_MODE_17                               = 0,
   parameter PINS_DATA_IN_MODE_18                               = 0,
   parameter PINS_DATA_IN_MODE_19                               = 0,
   parameter PINS_DATA_IN_MODE_20                               = 0,
   parameter PINS_DATA_IN_MODE_21                               = 0,
   parameter PINS_DATA_IN_MODE_22                               = 0,
   parameter PINS_DATA_IN_MODE_23                               = 0,
   parameter PINS_DATA_IN_MODE_24                               = 0,
   parameter PINS_DATA_IN_MODE_25                               = 0,
   parameter PINS_DATA_IN_MODE_26                               = 0,
   parameter PINS_DATA_IN_MODE_27                               = 0,
   parameter PINS_DATA_IN_MODE_28                               = 0,
   parameter PINS_DATA_IN_MODE_29                               = 0,
   parameter PINS_DATA_IN_MODE_30                               = 0,
   parameter PINS_DATA_IN_MODE_31                               = 0,
   parameter PINS_DATA_IN_MODE_32                               = 0,
   parameter PINS_DATA_IN_MODE_33                               = 0,
   parameter PINS_DATA_IN_MODE_34                               = 0,
   parameter PINS_DATA_IN_MODE_35                               = 0,
   parameter PINS_DATA_IN_MODE_36                               = 0,
   parameter PINS_DATA_IN_MODE_37                               = 0,
   parameter PINS_DATA_IN_MODE_38                               = 0,
   parameter PINS_DATA_IN_MODE_AUTOGEN_WCNT                     = 0,
   parameter PINS_C2L_DRIVEN_0                                  = 0,
   parameter PINS_C2L_DRIVEN_1                                  = 0,
   parameter PINS_C2L_DRIVEN_2                                  = 0,
   parameter PINS_C2L_DRIVEN_3                                  = 0,
   parameter PINS_C2L_DRIVEN_4                                  = 0,
   parameter PINS_C2L_DRIVEN_5                                  = 0,
   parameter PINS_C2L_DRIVEN_6                                  = 0,
   parameter PINS_C2L_DRIVEN_7                                  = 0,
   parameter PINS_C2L_DRIVEN_8                                  = 0,
   parameter PINS_C2L_DRIVEN_9                                  = 0,
   parameter PINS_C2L_DRIVEN_10                                 = 0,
   parameter PINS_C2L_DRIVEN_11                                 = 0,
   parameter PINS_C2L_DRIVEN_12                                 = 0,
   parameter PINS_C2L_DRIVEN_AUTOGEN_WCNT                       = 0,
   parameter PINS_DB_IN_BYPASS_0                                = 0,
   parameter PINS_DB_IN_BYPASS_1                                = 0,
   parameter PINS_DB_IN_BYPASS_2                                = 0,
   parameter PINS_DB_IN_BYPASS_3                                = 0,
   parameter PINS_DB_IN_BYPASS_4                                = 0,
   parameter PINS_DB_IN_BYPASS_5                                = 0,
   parameter PINS_DB_IN_BYPASS_6                                = 0,
   parameter PINS_DB_IN_BYPASS_7                                = 0,
   parameter PINS_DB_IN_BYPASS_8                                = 0,
   parameter PINS_DB_IN_BYPASS_9                                = 0,
   parameter PINS_DB_IN_BYPASS_10                               = 0,
   parameter PINS_DB_IN_BYPASS_11                               = 0,
   parameter PINS_DB_IN_BYPASS_12                               = 0,
   parameter PINS_DB_IN_BYPASS_AUTOGEN_WCNT                     = 0,
   parameter PINS_DB_OUT_BYPASS_0                               = 0,
   parameter PINS_DB_OUT_BYPASS_1                               = 0,
   parameter PINS_DB_OUT_BYPASS_2                               = 0,
   parameter PINS_DB_OUT_BYPASS_3                               = 0,
   parameter PINS_DB_OUT_BYPASS_4                               = 0,
   parameter PINS_DB_OUT_BYPASS_5                               = 0,
   parameter PINS_DB_OUT_BYPASS_6                               = 0,
   parameter PINS_DB_OUT_BYPASS_7                               = 0,
   parameter PINS_DB_OUT_BYPASS_8                               = 0,
   parameter PINS_DB_OUT_BYPASS_9                               = 0,
   parameter PINS_DB_OUT_BYPASS_10                              = 0,
   parameter PINS_DB_OUT_BYPASS_11                              = 0,
   parameter PINS_DB_OUT_BYPASS_12                              = 0,
   parameter PINS_DB_OUT_BYPASS_AUTOGEN_WCNT                    = 0,
   parameter PINS_DB_OE_BYPASS_0                                = 0,
   parameter PINS_DB_OE_BYPASS_1                                = 0,
   parameter PINS_DB_OE_BYPASS_2                                = 0,
   parameter PINS_DB_OE_BYPASS_3                                = 0,
   parameter PINS_DB_OE_BYPASS_4                                = 0,
   parameter PINS_DB_OE_BYPASS_5                                = 0,
   parameter PINS_DB_OE_BYPASS_6                                = 0,
   parameter PINS_DB_OE_BYPASS_7                                = 0,
   parameter PINS_DB_OE_BYPASS_8                                = 0,
   parameter PINS_DB_OE_BYPASS_9                                = 0,
   parameter PINS_DB_OE_BYPASS_10                               = 0,
   parameter PINS_DB_OE_BYPASS_11                               = 0,
   parameter PINS_DB_OE_BYPASS_12                               = 0,
   parameter PINS_DB_OE_BYPASS_AUTOGEN_WCNT                     = 0,
   parameter PINS_INVERT_WR_0                                   = 0,
   parameter PINS_INVERT_WR_1                                   = 0,
   parameter PINS_INVERT_WR_2                                   = 0,
   parameter PINS_INVERT_WR_3                                   = 0,
   parameter PINS_INVERT_WR_4                                   = 0,
   parameter PINS_INVERT_WR_5                                   = 0,
   parameter PINS_INVERT_WR_6                                   = 0,
   parameter PINS_INVERT_WR_7                                   = 0,
   parameter PINS_INVERT_WR_8                                   = 0,
   parameter PINS_INVERT_WR_9                                   = 0,
   parameter PINS_INVERT_WR_10                                  = 0,
   parameter PINS_INVERT_WR_11                                  = 0,
   parameter PINS_INVERT_WR_12                                  = 0,
   parameter PINS_INVERT_WR_AUTOGEN_WCNT                        = 0,
   parameter PINS_INVERT_OE_0                                   = 0,
   parameter PINS_INVERT_OE_1                                   = 0,
   parameter PINS_INVERT_OE_2                                   = 0,
   parameter PINS_INVERT_OE_3                                   = 0,
   parameter PINS_INVERT_OE_4                                   = 0,
   parameter PINS_INVERT_OE_5                                   = 0,
   parameter PINS_INVERT_OE_6                                   = 0,
   parameter PINS_INVERT_OE_7                                   = 0,
   parameter PINS_INVERT_OE_8                                   = 0,
   parameter PINS_INVERT_OE_9                                   = 0,
   parameter PINS_INVERT_OE_10                                  = 0,
   parameter PINS_INVERT_OE_11                                  = 0,
   parameter PINS_INVERT_OE_12                                  = 0,
   parameter PINS_INVERT_OE_AUTOGEN_WCNT                        = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_0                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_1                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_2                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_3                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_4                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_5                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_6                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_7                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_8                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_9                    = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_10                   = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_11                   = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_12                   = 0,
   parameter PINS_AC_HMC_DATA_OVERRIDE_ENA_AUTOGEN_WCNT         = 0,
   parameter PINS_OCT_MODE_0                                    = 0,
   parameter PINS_OCT_MODE_1                                    = 0,
   parameter PINS_OCT_MODE_2                                    = 0,
   parameter PINS_OCT_MODE_3                                    = 0,
   parameter PINS_OCT_MODE_4                                    = 0,
   parameter PINS_OCT_MODE_5                                    = 0,
   parameter PINS_OCT_MODE_6                                    = 0,
   parameter PINS_OCT_MODE_7                                    = 0,
   parameter PINS_OCT_MODE_8                                    = 0,
   parameter PINS_OCT_MODE_9                                    = 0,
   parameter PINS_OCT_MODE_10                                   = 0,
   parameter PINS_OCT_MODE_11                                   = 0,
   parameter PINS_OCT_MODE_12                                   = 0,
   parameter PINS_OCT_MODE_AUTOGEN_WCNT                         = 0,
   parameter PINS_GPIO_MODE_0                                   = 0,
   parameter PINS_GPIO_MODE_1                                   = 0,
   parameter PINS_GPIO_MODE_2                                   = 0,
   parameter PINS_GPIO_MODE_3                                   = 0,
   parameter PINS_GPIO_MODE_4                                   = 0,
   parameter PINS_GPIO_MODE_5                                   = 0,
   parameter PINS_GPIO_MODE_6                                   = 0,
   parameter PINS_GPIO_MODE_7                                   = 0,
   parameter PINS_GPIO_MODE_8                                   = 0,
   parameter PINS_GPIO_MODE_9                                   = 0,
   parameter PINS_GPIO_MODE_10                                  = 0,
   parameter PINS_GPIO_MODE_11                                  = 0,
   parameter PINS_GPIO_MODE_12                                  = 0,
   parameter PINS_GPIO_MODE_AUTOGEN_WCNT                        = 0,
   parameter UNUSED_MEM_PINS_PINLOC_0                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_1                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_2                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_3                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_4                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_5                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_6                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_7                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_8                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_9                           = 0,
   parameter UNUSED_MEM_PINS_PINLOC_10                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_11                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_12                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_13                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_14                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_15                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_16                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_17                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_18                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_19                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_20                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_21                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_22                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_23                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_24                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_25                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_26                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_27                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_28                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_29                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_30                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_31                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_32                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_33                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_34                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_35                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_36                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_37                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_38                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_39                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_40                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_41                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_42                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_43                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_44                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_45                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_46                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_47                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_48                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_49                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_50                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_51                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_52                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_53                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_54                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_55                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_56                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_57                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_58                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_59                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_60                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_61                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_62                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_63                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_64                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_65                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_66                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_67                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_68                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_69                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_70                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_71                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_72                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_73                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_74                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_75                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_76                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_77                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_78                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_79                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_80                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_81                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_82                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_83                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_84                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_85                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_86                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_87                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_88                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_89                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_90                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_91                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_92                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_93                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_94                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_95                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_96                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_97                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_98                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_99                          = 0,
   parameter UNUSED_MEM_PINS_PINLOC_100                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_101                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_102                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_103                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_104                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_105                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_106                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_107                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_108                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_109                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_110                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_111                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_112                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_113                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_114                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_115                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_116                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_117                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_118                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_119                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_120                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_121                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_122                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_123                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_124                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_125                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_126                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_127                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_128                         = 0,
   parameter UNUSED_MEM_PINS_PINLOC_AUTOGEN_WCNT                = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_0                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_1                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_2                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_3                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_4                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_5                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_6                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_7                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_8                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_9                         = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_10                        = 0,
   parameter UNUSED_DQS_BUSES_LANELOC_AUTOGEN_WCNT              = 0,
   parameter CENTER_TIDS_0                                      = 0,
   parameter CENTER_TIDS_1                                      = 0,
   parameter CENTER_TIDS_2                                      = 0,
   parameter CENTER_TIDS_AUTOGEN_WCNT                           = 0,
   parameter HMC_TIDS_0                                         = 0,
   parameter HMC_TIDS_1                                         = 0,
   parameter HMC_TIDS_2                                         = 0,
   parameter HMC_TIDS_AUTOGEN_WCNT                              = 0,
   parameter LANE_TIDS_0                                        = 0,
   parameter LANE_TIDS_1                                        = 0,
   parameter LANE_TIDS_2                                        = 0,
   parameter LANE_TIDS_3                                        = 0,
   parameter LANE_TIDS_4                                        = 0,
   parameter LANE_TIDS_5                                        = 0,
   parameter LANE_TIDS_6                                        = 0,
   parameter LANE_TIDS_7                                        = 0,
   parameter LANE_TIDS_8                                        = 0,
   parameter LANE_TIDS_9                                        = 0,
   parameter LANE_TIDS_AUTOGEN_WCNT                             = 0,
   parameter PREAMBLE_MODE                                      = "",
   parameter DBI_WR_ENABLE                                      = "",
   parameter DBI_RD_ENABLE                                      = "",
   parameter CRC_EN                                             = "",
   parameter SWAP_DQS_A_B                                       = "",
   parameter DQS_PACK_MODE                                      = "",
   parameter OCT_SIZE                                           = 0,
   parameter DBC_WB_RESERVED_ENTRY                              = 0,
   parameter DLL_MODE                                           = "",
   parameter DLL_CODEWORD                                       = 0,
   parameter ABPHY_WRITE_PROTOCOL                               = 0,
   parameter PHY_USERMODE_OCT                                   = 0,
   parameter PHY_PERIODIC_OCT_RECAL                             = 0,
   parameter PHY_HAS_DCC                                        = 0,
   parameter PRI_HMC_CFG_ENABLE_ECC                             = "",
   parameter PRI_HMC_CFG_REORDER_DATA                           = "",
   parameter PRI_HMC_CFG_REORDER_READ                           = "",
   parameter PRI_HMC_CFG_REORDER_RDATA                          = "",
   parameter PRI_HMC_CFG_STARVE_LIMIT                           = 0,
   parameter PRI_HMC_CFG_DQS_TRACKING_EN                        = "",
   parameter PRI_HMC_CFG_ARBITER_TYPE                           = "",
   parameter PRI_HMC_CFG_OPEN_PAGE_EN                           = "",
   parameter PRI_HMC_CFG_GEAR_DOWN_EN                           = "",
   parameter PRI_HMC_CFG_RLD3_MULTIBANK_MODE                    = "",
   parameter PRI_HMC_CFG_PING_PONG_MODE                         = "",
   parameter PRI_HMC_CFG_SLOT_ROTATE_EN                         = 0,
   parameter PRI_HMC_CFG_SLOT_OFFSET                            = 0,
   parameter PRI_HMC_CFG_COL_CMD_SLOT                           = 0,
   parameter PRI_HMC_CFG_ROW_CMD_SLOT                           = 0,
   parameter PRI_HMC_CFG_ENABLE_RC                              = "",
   parameter PRI_HMC_CFG_CS_TO_CHIP_MAPPING                     = 0,
   parameter PRI_HMC_CFG_RB_RESERVED_ENTRY                      = 0,
   parameter PRI_HMC_CFG_WB_RESERVED_ENTRY                      = 0,
   parameter PRI_HMC_CFG_TCL                                    = 0,
   parameter PRI_HMC_CFG_POWER_SAVING_EXIT_CYC                  = 0,
   parameter PRI_HMC_CFG_MEM_CLK_DISABLE_ENTRY_CYC              = 0,
   parameter PRI_HMC_CFG_WRITE_ODT_CHIP                         = 0,
   parameter PRI_HMC_CFG_READ_ODT_CHIP                          = 0,
   parameter PRI_HMC_CFG_WR_ODT_ON                              = 0,
   parameter PRI_HMC_CFG_RD_ODT_ON                              = 0,
   parameter PRI_HMC_CFG_WR_ODT_PERIOD                          = 0,
   parameter PRI_HMC_CFG_RD_ODT_PERIOD                          = 0,
   parameter PRI_HMC_CFG_RLD3_REFRESH_SEQ0                      = 0,
   parameter PRI_HMC_CFG_RLD3_REFRESH_SEQ1                      = 0,
   parameter PRI_HMC_CFG_RLD3_REFRESH_SEQ2                      = 0,
   parameter PRI_HMC_CFG_RLD3_REFRESH_SEQ3                      = 0,
   parameter PRI_HMC_CFG_SRF_ZQCAL_DISABLE                      = "",
   parameter PRI_HMC_CFG_MPS_ZQCAL_DISABLE                      = "",
   parameter PRI_HMC_CFG_MPS_DQSTRK_DISABLE                     = "",
   parameter PRI_HMC_CFG_SHORT_DQSTRK_CTRL_EN                   = "",
   parameter PRI_HMC_CFG_PERIOD_DQSTRK_CTRL_EN                  = "",
   parameter PRI_HMC_CFG_PERIOD_DQSTRK_INTERVAL                 = 0,
   parameter PRI_HMC_CFG_DQSTRK_TO_VALID_LAST                   = 0,
   parameter PRI_HMC_CFG_DQSTRK_TO_VALID                        = 0,
   parameter PRI_HMC_CFG_RFSH_WARN_THRESHOLD                    = 0,
   parameter PRI_HMC_CFG_SB_CG_DISABLE                          = "",
   parameter PRI_HMC_CFG_USER_RFSH_EN                           = "",
   parameter PRI_HMC_CFG_SRF_AUTOEXIT_EN                        = "",
   parameter PRI_HMC_CFG_SRF_ENTRY_EXIT_BLOCK                   = "",
   parameter PRI_HMC_CFG_SB_DDR4_MR3                            = 0,
   parameter PRI_HMC_CFG_SB_DDR4_MR4                            = 0,
   parameter PRI_HMC_CFG_SB_DDR4_MR5                            = 0,
   parameter PRI_HMC_CFG_DDR4_MPS_ADDR_MIRROR                   = 0,
   parameter PRI_HMC_CFG_MEM_IF_COLADDR_WIDTH                   = "",
   parameter PRI_HMC_CFG_MEM_IF_ROWADDR_WIDTH                   = "",
   parameter PRI_HMC_CFG_MEM_IF_BANKADDR_WIDTH                  = "",
   parameter PRI_HMC_CFG_MEM_IF_BGADDR_WIDTH                    = "",
   parameter PRI_HMC_CFG_LOCAL_IF_CS_WIDTH                      = "",
   parameter PRI_HMC_CFG_ADDR_ORDER                             = "",
   parameter PRI_HMC_CFG_ACT_TO_RDWR                            = 0,
   parameter PRI_HMC_CFG_ACT_TO_PCH                             = 0,
   parameter PRI_HMC_CFG_ACT_TO_ACT                             = 0,
   parameter PRI_HMC_CFG_ACT_TO_ACT_DIFF_BANK                   = 0,
   parameter PRI_HMC_CFG_ACT_TO_ACT_DIFF_BG                     = 0,
   parameter PRI_HMC_CFG_RD_TO_RD                               = 0,
   parameter PRI_HMC_CFG_RD_TO_RD_DIFF_CHIP                     = 0,
   parameter PRI_HMC_CFG_RD_TO_RD_DIFF_BG                       = 0,
   parameter PRI_HMC_CFG_RD_TO_WR                               = 0,
   parameter PRI_HMC_CFG_RD_TO_WR_DIFF_CHIP                     = 0,
   parameter PRI_HMC_CFG_RD_TO_WR_DIFF_BG                       = 0,
   parameter PRI_HMC_CFG_RD_TO_PCH                              = 0,
   parameter PRI_HMC_CFG_RD_AP_TO_VALID                         = 0,
   parameter PRI_HMC_CFG_WR_TO_WR                               = 0,
   parameter PRI_HMC_CFG_WR_TO_WR_DIFF_CHIP                     = 0,
   parameter PRI_HMC_CFG_WR_TO_WR_DIFF_BG                       = 0,
   parameter PRI_HMC_CFG_WR_TO_RD                               = 0,
   parameter PRI_HMC_CFG_WR_TO_RD_DIFF_CHIP                     = 0,
   parameter PRI_HMC_CFG_WR_TO_RD_DIFF_BG                       = 0,
   parameter PRI_HMC_CFG_WR_TO_PCH                              = 0,
   parameter PRI_HMC_CFG_WR_AP_TO_VALID                         = 0,
   parameter PRI_HMC_CFG_PCH_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_PCH_ALL_TO_VALID                       = 0,
   parameter PRI_HMC_CFG_ARF_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_PDN_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_SRF_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_SRF_TO_ZQ_CAL                          = 0,
   parameter PRI_HMC_CFG_ARF_PERIOD                             = 0,
   parameter PRI_HMC_CFG_PDN_PERIOD                             = 0,
   parameter PRI_HMC_CFG_ZQCL_TO_VALID                          = 0,
   parameter PRI_HMC_CFG_ZQCS_TO_VALID                          = 0,
   parameter PRI_HMC_CFG_MRS_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_MPS_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_MRR_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_MPR_TO_VALID                           = 0,
   parameter PRI_HMC_CFG_MPS_EXIT_CS_TO_CKE                     = 0,
   parameter PRI_HMC_CFG_MPS_EXIT_CKE_TO_CS                     = 0,
   parameter PRI_HMC_CFG_RLD3_MULTIBANK_REF_DELAY               = 0,
   parameter PRI_HMC_CFG_MMR_CMD_TO_VALID                       = 0,
   parameter PRI_HMC_CFG_4_ACT_TO_ACT                           = 0,
   parameter PRI_HMC_CFG_16_ACT_TO_ACT                          = 0,
   parameter SEC_HMC_CFG_ENABLE_ECC                             = "",
   parameter SEC_HMC_CFG_REORDER_DATA                           = "",
   parameter SEC_HMC_CFG_REORDER_READ                           = "",
   parameter SEC_HMC_CFG_REORDER_RDATA                          = "",
   parameter SEC_HMC_CFG_STARVE_LIMIT                           = 0,
   parameter SEC_HMC_CFG_DQS_TRACKING_EN                        = "",
   parameter SEC_HMC_CFG_ARBITER_TYPE                           = "",
   parameter SEC_HMC_CFG_OPEN_PAGE_EN                           = "",
   parameter SEC_HMC_CFG_GEAR_DOWN_EN                           = "",
   parameter SEC_HMC_CFG_RLD3_MULTIBANK_MODE                    = "",
   parameter SEC_HMC_CFG_PING_PONG_MODE                         = "",
   parameter SEC_HMC_CFG_SLOT_ROTATE_EN                         = 0,
   parameter SEC_HMC_CFG_SLOT_OFFSET                            = 0,
   parameter SEC_HMC_CFG_COL_CMD_SLOT                           = 0,
   parameter SEC_HMC_CFG_ROW_CMD_SLOT                           = 0,
   parameter SEC_HMC_CFG_ENABLE_RC                              = "",
   parameter SEC_HMC_CFG_CS_TO_CHIP_MAPPING                     = 0,
   parameter SEC_HMC_CFG_RB_RESERVED_ENTRY                      = 0,
   parameter SEC_HMC_CFG_WB_RESERVED_ENTRY                      = 0,
   parameter SEC_HMC_CFG_TCL                                    = 0,
   parameter SEC_HMC_CFG_POWER_SAVING_EXIT_CYC                  = 0,
   parameter SEC_HMC_CFG_MEM_CLK_DISABLE_ENTRY_CYC              = 0,
   parameter SEC_HMC_CFG_WRITE_ODT_CHIP                         = 0,
   parameter SEC_HMC_CFG_READ_ODT_CHIP                          = 0,
   parameter SEC_HMC_CFG_WR_ODT_ON                              = 0,
   parameter SEC_HMC_CFG_RD_ODT_ON                              = 0,
   parameter SEC_HMC_CFG_WR_ODT_PERIOD                          = 0,
   parameter SEC_HMC_CFG_RD_ODT_PERIOD                          = 0,
   parameter SEC_HMC_CFG_RLD3_REFRESH_SEQ0                      = 0,
   parameter SEC_HMC_CFG_RLD3_REFRESH_SEQ1                      = 0,
   parameter SEC_HMC_CFG_RLD3_REFRESH_SEQ2                      = 0,
   parameter SEC_HMC_CFG_RLD3_REFRESH_SEQ3                      = 0,
   parameter SEC_HMC_CFG_SRF_ZQCAL_DISABLE                      = "",
   parameter SEC_HMC_CFG_MPS_ZQCAL_DISABLE                      = "",
   parameter SEC_HMC_CFG_MPS_DQSTRK_DISABLE                     = "",
   parameter SEC_HMC_CFG_SHORT_DQSTRK_CTRL_EN                   = "",
   parameter SEC_HMC_CFG_PERIOD_DQSTRK_CTRL_EN                  = "",
   parameter SEC_HMC_CFG_PERIOD_DQSTRK_INTERVAL                 = 0,
   parameter SEC_HMC_CFG_DQSTRK_TO_VALID_LAST                   = 0,
   parameter SEC_HMC_CFG_DQSTRK_TO_VALID                        = 0,
   parameter SEC_HMC_CFG_RFSH_WARN_THRESHOLD                    = 0,
   parameter SEC_HMC_CFG_SB_CG_DISABLE                          = "",
   parameter SEC_HMC_CFG_USER_RFSH_EN                           = "",
   parameter SEC_HMC_CFG_SRF_AUTOEXIT_EN                        = "",
   parameter SEC_HMC_CFG_SRF_ENTRY_EXIT_BLOCK                   = "",
   parameter SEC_HMC_CFG_SB_DDR4_MR3                            = 0,
   parameter SEC_HMC_CFG_SB_DDR4_MR4                            = 0,
   parameter SEC_HMC_CFG_SB_DDR4_MR5                            = 0,
   parameter SEC_HMC_CFG_DDR4_MPS_ADDR_MIRROR                   = 0,
   parameter SEC_HMC_CFG_MEM_IF_COLADDR_WIDTH                   = "",
   parameter SEC_HMC_CFG_MEM_IF_ROWADDR_WIDTH                   = "",
   parameter SEC_HMC_CFG_MEM_IF_BANKADDR_WIDTH                  = "",
   parameter SEC_HMC_CFG_MEM_IF_BGADDR_WIDTH                    = "",
   parameter SEC_HMC_CFG_LOCAL_IF_CS_WIDTH                      = "",
   parameter SEC_HMC_CFG_ADDR_ORDER                             = "",
   parameter SEC_HMC_CFG_ACT_TO_RDWR                            = 0,
   parameter SEC_HMC_CFG_ACT_TO_PCH                             = 0,
   parameter SEC_HMC_CFG_ACT_TO_ACT                             = 0,
   parameter SEC_HMC_CFG_ACT_TO_ACT_DIFF_BANK                   = 0,
   parameter SEC_HMC_CFG_ACT_TO_ACT_DIFF_BG                     = 0,
   parameter SEC_HMC_CFG_RD_TO_RD                               = 0,
   parameter SEC_HMC_CFG_RD_TO_RD_DIFF_CHIP                     = 0,
   parameter SEC_HMC_CFG_RD_TO_RD_DIFF_BG                       = 0,
   parameter SEC_HMC_CFG_RD_TO_WR                               = 0,
   parameter SEC_HMC_CFG_RD_TO_WR_DIFF_CHIP                     = 0,
   parameter SEC_HMC_CFG_RD_TO_WR_DIFF_BG                       = 0,
   parameter SEC_HMC_CFG_RD_TO_PCH                              = 0,
   parameter SEC_HMC_CFG_RD_AP_TO_VALID                         = 0,
   parameter SEC_HMC_CFG_WR_TO_WR                               = 0,
   parameter SEC_HMC_CFG_WR_TO_WR_DIFF_CHIP                     = 0,
   parameter SEC_HMC_CFG_WR_TO_WR_DIFF_BG                       = 0,
   parameter SEC_HMC_CFG_WR_TO_RD                               = 0,
   parameter SEC_HMC_CFG_WR_TO_RD_DIFF_CHIP                     = 0,
   parameter SEC_HMC_CFG_WR_TO_RD_DIFF_BG                       = 0,
   parameter SEC_HMC_CFG_WR_TO_PCH                              = 0,
   parameter SEC_HMC_CFG_WR_AP_TO_VALID                         = 0,
   parameter SEC_HMC_CFG_PCH_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_PCH_ALL_TO_VALID                       = 0,
   parameter SEC_HMC_CFG_ARF_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_PDN_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_SRF_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_SRF_TO_ZQ_CAL                          = 0,
   parameter SEC_HMC_CFG_ARF_PERIOD                             = 0,
   parameter SEC_HMC_CFG_PDN_PERIOD                             = 0,
   parameter SEC_HMC_CFG_ZQCL_TO_VALID                          = 0,
   parameter SEC_HMC_CFG_ZQCS_TO_VALID                          = 0,
   parameter SEC_HMC_CFG_MRS_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_MPS_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_MRR_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_MPR_TO_VALID                           = 0,
   parameter SEC_HMC_CFG_MPS_EXIT_CS_TO_CKE                     = 0,
   parameter SEC_HMC_CFG_MPS_EXIT_CKE_TO_CS                     = 0,
   parameter SEC_HMC_CFG_RLD3_MULTIBANK_REF_DELAY               = 0,
   parameter SEC_HMC_CFG_MMR_CMD_TO_VALID                       = 0,
   parameter SEC_HMC_CFG_4_ACT_TO_ACT                           = 0,
   parameter SEC_HMC_CFG_16_ACT_TO_ACT                          = 0,
   parameter PINS_PER_LANE                                      = 0,
   parameter LANES_PER_TILE                                     = 0,
   parameter OCT_CONTROL_WIDTH                                  = 0,
   parameter PORT_MEM_CK_WIDTH                                  = 0,
   parameter PORT_MEM_CK_PINLOC_0                               = 0,
   parameter PORT_MEM_CK_PINLOC_1                               = 0,
   parameter PORT_MEM_CK_PINLOC_2                               = 0,
   parameter PORT_MEM_CK_PINLOC_3                               = 0,
   parameter PORT_MEM_CK_PINLOC_4                               = 0,
   parameter PORT_MEM_CK_PINLOC_5                               = 0,
   parameter PORT_MEM_CK_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_CK_N_WIDTH                                = 0,
   parameter PORT_MEM_CK_N_PINLOC_0                             = 0,
   parameter PORT_MEM_CK_N_PINLOC_1                             = 0,
   parameter PORT_MEM_CK_N_PINLOC_2                             = 0,
   parameter PORT_MEM_CK_N_PINLOC_3                             = 0,
   parameter PORT_MEM_CK_N_PINLOC_4                             = 0,
   parameter PORT_MEM_CK_N_PINLOC_5                             = 0,
   parameter PORT_MEM_CK_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_DK_WIDTH                                  = 0,
   parameter PORT_MEM_DK_PINLOC_0                               = 0,
   parameter PORT_MEM_DK_PINLOC_1                               = 0,
   parameter PORT_MEM_DK_PINLOC_2                               = 0,
   parameter PORT_MEM_DK_PINLOC_3                               = 0,
   parameter PORT_MEM_DK_PINLOC_4                               = 0,
   parameter PORT_MEM_DK_PINLOC_5                               = 0,
   parameter PORT_MEM_DK_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_DK_N_WIDTH                                = 0,
   parameter PORT_MEM_DK_N_PINLOC_0                             = 0,
   parameter PORT_MEM_DK_N_PINLOC_1                             = 0,
   parameter PORT_MEM_DK_N_PINLOC_2                             = 0,
   parameter PORT_MEM_DK_N_PINLOC_3                             = 0,
   parameter PORT_MEM_DK_N_PINLOC_4                             = 0,
   parameter PORT_MEM_DK_N_PINLOC_5                             = 0,
   parameter PORT_MEM_DK_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_DKA_WIDTH                                 = 0,
   parameter PORT_MEM_DKA_PINLOC_0                              = 0,
   parameter PORT_MEM_DKA_PINLOC_1                              = 0,
   parameter PORT_MEM_DKA_PINLOC_2                              = 0,
   parameter PORT_MEM_DKA_PINLOC_3                              = 0,
   parameter PORT_MEM_DKA_PINLOC_4                              = 0,
   parameter PORT_MEM_DKA_PINLOC_5                              = 0,
   parameter PORT_MEM_DKA_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_DKA_N_WIDTH                               = 0,
   parameter PORT_MEM_DKA_N_PINLOC_0                            = 0,
   parameter PORT_MEM_DKA_N_PINLOC_1                            = 0,
   parameter PORT_MEM_DKA_N_PINLOC_2                            = 0,
   parameter PORT_MEM_DKA_N_PINLOC_3                            = 0,
   parameter PORT_MEM_DKA_N_PINLOC_4                            = 0,
   parameter PORT_MEM_DKA_N_PINLOC_5                            = 0,
   parameter PORT_MEM_DKA_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_DKB_WIDTH                                 = 0,
   parameter PORT_MEM_DKB_PINLOC_0                              = 0,
   parameter PORT_MEM_DKB_PINLOC_1                              = 0,
   parameter PORT_MEM_DKB_PINLOC_2                              = 0,
   parameter PORT_MEM_DKB_PINLOC_3                              = 0,
   parameter PORT_MEM_DKB_PINLOC_4                              = 0,
   parameter PORT_MEM_DKB_PINLOC_5                              = 0,
   parameter PORT_MEM_DKB_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_DKB_N_WIDTH                               = 0,
   parameter PORT_MEM_DKB_N_PINLOC_0                            = 0,
   parameter PORT_MEM_DKB_N_PINLOC_1                            = 0,
   parameter PORT_MEM_DKB_N_PINLOC_2                            = 0,
   parameter PORT_MEM_DKB_N_PINLOC_3                            = 0,
   parameter PORT_MEM_DKB_N_PINLOC_4                            = 0,
   parameter PORT_MEM_DKB_N_PINLOC_5                            = 0,
   parameter PORT_MEM_DKB_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_K_WIDTH                                   = 0,
   parameter PORT_MEM_K_PINLOC_0                                = 0,
   parameter PORT_MEM_K_PINLOC_1                                = 0,
   parameter PORT_MEM_K_PINLOC_2                                = 0,
   parameter PORT_MEM_K_PINLOC_3                                = 0,
   parameter PORT_MEM_K_PINLOC_4                                = 0,
   parameter PORT_MEM_K_PINLOC_5                                = 0,
   parameter PORT_MEM_K_PINLOC_AUTOGEN_WCNT                     = 0,
   parameter PORT_MEM_K_N_WIDTH                                 = 0,
   parameter PORT_MEM_K_N_PINLOC_0                              = 0,
   parameter PORT_MEM_K_N_PINLOC_1                              = 0,
   parameter PORT_MEM_K_N_PINLOC_2                              = 0,
   parameter PORT_MEM_K_N_PINLOC_3                              = 0,
   parameter PORT_MEM_K_N_PINLOC_4                              = 0,
   parameter PORT_MEM_K_N_PINLOC_5                              = 0,
   parameter PORT_MEM_K_N_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_A_WIDTH                                   = 0,
   parameter PORT_MEM_A_PINLOC_0                                = 0,
   parameter PORT_MEM_A_PINLOC_1                                = 0,
   parameter PORT_MEM_A_PINLOC_2                                = 0,
   parameter PORT_MEM_A_PINLOC_3                                = 0,
   parameter PORT_MEM_A_PINLOC_4                                = 0,
   parameter PORT_MEM_A_PINLOC_5                                = 0,
   parameter PORT_MEM_A_PINLOC_6                                = 0,
   parameter PORT_MEM_A_PINLOC_7                                = 0,
   parameter PORT_MEM_A_PINLOC_8                                = 0,
   parameter PORT_MEM_A_PINLOC_9                                = 0,
   parameter PORT_MEM_A_PINLOC_10                               = 0,
   parameter PORT_MEM_A_PINLOC_11                               = 0,
   parameter PORT_MEM_A_PINLOC_12                               = 0,
   parameter PORT_MEM_A_PINLOC_13                               = 0,
   parameter PORT_MEM_A_PINLOC_14                               = 0,
   parameter PORT_MEM_A_PINLOC_15                               = 0,
   parameter PORT_MEM_A_PINLOC_16                               = 0,
   parameter PORT_MEM_A_PINLOC_AUTOGEN_WCNT                     = 0,
   parameter PORT_MEM_BA_WIDTH                                  = 0,
   parameter PORT_MEM_BA_PINLOC_0                               = 0,
   parameter PORT_MEM_BA_PINLOC_1                               = 0,
   parameter PORT_MEM_BA_PINLOC_2                               = 0,
   parameter PORT_MEM_BA_PINLOC_3                               = 0,
   parameter PORT_MEM_BA_PINLOC_4                               = 0,
   parameter PORT_MEM_BA_PINLOC_5                               = 0,
   parameter PORT_MEM_BA_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_BG_WIDTH                                  = 0,
   parameter PORT_MEM_BG_PINLOC_0                               = 0,
   parameter PORT_MEM_BG_PINLOC_1                               = 0,
   parameter PORT_MEM_BG_PINLOC_2                               = 0,
   parameter PORT_MEM_BG_PINLOC_3                               = 0,
   parameter PORT_MEM_BG_PINLOC_4                               = 0,
   parameter PORT_MEM_BG_PINLOC_5                               = 0,
   parameter PORT_MEM_BG_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_C_WIDTH                                   = 0,
   parameter PORT_MEM_C_PINLOC_0                                = 0,
   parameter PORT_MEM_C_PINLOC_1                                = 0,
   parameter PORT_MEM_C_PINLOC_2                                = 0,
   parameter PORT_MEM_C_PINLOC_3                                = 0,
   parameter PORT_MEM_C_PINLOC_4                                = 0,
   parameter PORT_MEM_C_PINLOC_5                                = 0,
   parameter PORT_MEM_C_PINLOC_AUTOGEN_WCNT                     = 0,
   parameter PORT_MEM_CKE_WIDTH                                 = 0,
   parameter PORT_MEM_CKE_PINLOC_0                              = 0,
   parameter PORT_MEM_CKE_PINLOC_1                              = 0,
   parameter PORT_MEM_CKE_PINLOC_2                              = 0,
   parameter PORT_MEM_CKE_PINLOC_3                              = 0,
   parameter PORT_MEM_CKE_PINLOC_4                              = 0,
   parameter PORT_MEM_CKE_PINLOC_5                              = 0,
   parameter PORT_MEM_CKE_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_CS_N_WIDTH                                = 0,
   parameter PORT_MEM_CS_N_PINLOC_0                             = 0,
   parameter PORT_MEM_CS_N_PINLOC_1                             = 0,
   parameter PORT_MEM_CS_N_PINLOC_2                             = 0,
   parameter PORT_MEM_CS_N_PINLOC_3                             = 0,
   parameter PORT_MEM_CS_N_PINLOC_4                             = 0,
   parameter PORT_MEM_CS_N_PINLOC_5                             = 0,
   parameter PORT_MEM_CS_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_RM_WIDTH                                  = 0,
   parameter PORT_MEM_RM_PINLOC_0                               = 0,
   parameter PORT_MEM_RM_PINLOC_1                               = 0,
   parameter PORT_MEM_RM_PINLOC_2                               = 0,
   parameter PORT_MEM_RM_PINLOC_3                               = 0,
   parameter PORT_MEM_RM_PINLOC_4                               = 0,
   parameter PORT_MEM_RM_PINLOC_5                               = 0,
   parameter PORT_MEM_RM_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_ODT_WIDTH                                 = 0,
   parameter PORT_MEM_ODT_PINLOC_0                              = 0,
   parameter PORT_MEM_ODT_PINLOC_1                              = 0,
   parameter PORT_MEM_ODT_PINLOC_2                              = 0,
   parameter PORT_MEM_ODT_PINLOC_3                              = 0,
   parameter PORT_MEM_ODT_PINLOC_4                              = 0,
   parameter PORT_MEM_ODT_PINLOC_5                              = 0,
   parameter PORT_MEM_ODT_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_RAS_N_WIDTH                               = 0,
   parameter PORT_MEM_RAS_N_PINLOC_0                            = 0,
   parameter PORT_MEM_RAS_N_PINLOC_1                            = 0,
   parameter PORT_MEM_RAS_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_CAS_N_WIDTH                               = 0,
   parameter PORT_MEM_CAS_N_PINLOC_0                            = 0,
   parameter PORT_MEM_CAS_N_PINLOC_1                            = 0,
   parameter PORT_MEM_CAS_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_WE_N_WIDTH                                = 0,
   parameter PORT_MEM_WE_N_PINLOC_0                             = 0,
   parameter PORT_MEM_WE_N_PINLOC_1                             = 0,
   parameter PORT_MEM_WE_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_RESET_N_WIDTH                             = 0,
   parameter PORT_MEM_RESET_N_PINLOC_0                          = 0,
   parameter PORT_MEM_RESET_N_PINLOC_1                          = 0,
   parameter PORT_MEM_RESET_N_PINLOC_AUTOGEN_WCNT               = 0,
   parameter PORT_MEM_ACT_N_WIDTH                               = 0,
   parameter PORT_MEM_ACT_N_PINLOC_0                            = 0,
   parameter PORT_MEM_ACT_N_PINLOC_1                            = 0,
   parameter PORT_MEM_ACT_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_PAR_WIDTH                                 = 0,
   parameter PORT_MEM_PAR_PINLOC_0                              = 0,
   parameter PORT_MEM_PAR_PINLOC_1                              = 0,
   parameter PORT_MEM_PAR_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_CA_WIDTH                                  = 0,
   parameter PORT_MEM_CA_PINLOC_0                               = 0,
   parameter PORT_MEM_CA_PINLOC_1                               = 0,
   parameter PORT_MEM_CA_PINLOC_2                               = 0,
   parameter PORT_MEM_CA_PINLOC_3                               = 0,
   parameter PORT_MEM_CA_PINLOC_4                               = 0,
   parameter PORT_MEM_CA_PINLOC_5                               = 0,
   parameter PORT_MEM_CA_PINLOC_6                               = 0,
   parameter PORT_MEM_CA_PINLOC_7                               = 0,
   parameter PORT_MEM_CA_PINLOC_8                               = 0,
   parameter PORT_MEM_CA_PINLOC_9                               = 0,
   parameter PORT_MEM_CA_PINLOC_10                              = 0,
   parameter PORT_MEM_CA_PINLOC_11                              = 0,
   parameter PORT_MEM_CA_PINLOC_12                              = 0,
   parameter PORT_MEM_CA_PINLOC_13                              = 0,
   parameter PORT_MEM_CA_PINLOC_14                              = 0,
   parameter PORT_MEM_CA_PINLOC_15                              = 0,
   parameter PORT_MEM_CA_PINLOC_16                              = 0,
   parameter PORT_MEM_CA_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_REF_N_WIDTH                               = 0,
   parameter PORT_MEM_REF_N_PINLOC_0                            = 0,
   parameter PORT_MEM_REF_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_WPS_N_WIDTH                               = 0,
   parameter PORT_MEM_WPS_N_PINLOC_0                            = 0,
   parameter PORT_MEM_WPS_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_RPS_N_WIDTH                               = 0,
   parameter PORT_MEM_RPS_N_PINLOC_0                            = 0,
   parameter PORT_MEM_RPS_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_DOFF_N_WIDTH                              = 0,
   parameter PORT_MEM_DOFF_N_PINLOC_0                           = 0,
   parameter PORT_MEM_DOFF_N_PINLOC_AUTOGEN_WCNT                = 0,
   parameter PORT_MEM_LDA_N_WIDTH                               = 0,
   parameter PORT_MEM_LDA_N_PINLOC_0                            = 0,
   parameter PORT_MEM_LDA_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_LDB_N_WIDTH                               = 0,
   parameter PORT_MEM_LDB_N_PINLOC_0                            = 0,
   parameter PORT_MEM_LDB_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_RWA_N_WIDTH                               = 0,
   parameter PORT_MEM_RWA_N_PINLOC_0                            = 0,
   parameter PORT_MEM_RWA_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_RWB_N_WIDTH                               = 0,
   parameter PORT_MEM_RWB_N_PINLOC_0                            = 0,
   parameter PORT_MEM_RWB_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_LBK0_N_WIDTH                              = 0,
   parameter PORT_MEM_LBK0_N_PINLOC_0                           = 0,
   parameter PORT_MEM_LBK0_N_PINLOC_AUTOGEN_WCNT                = 0,
   parameter PORT_MEM_LBK1_N_WIDTH                              = 0,
   parameter PORT_MEM_LBK1_N_PINLOC_0                           = 0,
   parameter PORT_MEM_LBK1_N_PINLOC_AUTOGEN_WCNT                = 0,
   parameter PORT_MEM_CFG_N_WIDTH                               = 0,
   parameter PORT_MEM_CFG_N_PINLOC_0                            = 0,
   parameter PORT_MEM_CFG_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_AP_WIDTH                                  = 0,
   parameter PORT_MEM_AP_PINLOC_0                               = 0,
   parameter PORT_MEM_AP_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_AINV_WIDTH                                = 0,
   parameter PORT_MEM_AINV_PINLOC_0                             = 0,
   parameter PORT_MEM_AINV_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_DM_WIDTH                                  = 0,
   parameter PORT_MEM_DM_PINLOC_0                               = 0,
   parameter PORT_MEM_DM_PINLOC_1                               = 0,
   parameter PORT_MEM_DM_PINLOC_2                               = 0,
   parameter PORT_MEM_DM_PINLOC_3                               = 0,
   parameter PORT_MEM_DM_PINLOC_4                               = 0,
   parameter PORT_MEM_DM_PINLOC_5                               = 0,
   parameter PORT_MEM_DM_PINLOC_6                               = 0,
   parameter PORT_MEM_DM_PINLOC_7                               = 0,
   parameter PORT_MEM_DM_PINLOC_8                               = 0,
   parameter PORT_MEM_DM_PINLOC_9                               = 0,
   parameter PORT_MEM_DM_PINLOC_10                              = 0,
   parameter PORT_MEM_DM_PINLOC_11                              = 0,
   parameter PORT_MEM_DM_PINLOC_12                              = 0,
   parameter PORT_MEM_DM_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_BWS_N_WIDTH                               = 0,
   parameter PORT_MEM_BWS_N_PINLOC_0                            = 0,
   parameter PORT_MEM_BWS_N_PINLOC_1                            = 0,
   parameter PORT_MEM_BWS_N_PINLOC_2                            = 0,
   parameter PORT_MEM_BWS_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_D_WIDTH                                   = 0,
   parameter PORT_MEM_D_PINLOC_0                                = 0,
   parameter PORT_MEM_D_PINLOC_1                                = 0,
   parameter PORT_MEM_D_PINLOC_2                                = 0,
   parameter PORT_MEM_D_PINLOC_3                                = 0,
   parameter PORT_MEM_D_PINLOC_4                                = 0,
   parameter PORT_MEM_D_PINLOC_5                                = 0,
   parameter PORT_MEM_D_PINLOC_6                                = 0,
   parameter PORT_MEM_D_PINLOC_7                                = 0,
   parameter PORT_MEM_D_PINLOC_8                                = 0,
   parameter PORT_MEM_D_PINLOC_9                                = 0,
   parameter PORT_MEM_D_PINLOC_10                               = 0,
   parameter PORT_MEM_D_PINLOC_11                               = 0,
   parameter PORT_MEM_D_PINLOC_12                               = 0,
   parameter PORT_MEM_D_PINLOC_13                               = 0,
   parameter PORT_MEM_D_PINLOC_14                               = 0,
   parameter PORT_MEM_D_PINLOC_15                               = 0,
   parameter PORT_MEM_D_PINLOC_16                               = 0,
   parameter PORT_MEM_D_PINLOC_17                               = 0,
   parameter PORT_MEM_D_PINLOC_18                               = 0,
   parameter PORT_MEM_D_PINLOC_19                               = 0,
   parameter PORT_MEM_D_PINLOC_20                               = 0,
   parameter PORT_MEM_D_PINLOC_21                               = 0,
   parameter PORT_MEM_D_PINLOC_22                               = 0,
   parameter PORT_MEM_D_PINLOC_23                               = 0,
   parameter PORT_MEM_D_PINLOC_24                               = 0,
   parameter PORT_MEM_D_PINLOC_25                               = 0,
   parameter PORT_MEM_D_PINLOC_26                               = 0,
   parameter PORT_MEM_D_PINLOC_27                               = 0,
   parameter PORT_MEM_D_PINLOC_28                               = 0,
   parameter PORT_MEM_D_PINLOC_29                               = 0,
   parameter PORT_MEM_D_PINLOC_30                               = 0,
   parameter PORT_MEM_D_PINLOC_31                               = 0,
   parameter PORT_MEM_D_PINLOC_32                               = 0,
   parameter PORT_MEM_D_PINLOC_33                               = 0,
   parameter PORT_MEM_D_PINLOC_34                               = 0,
   parameter PORT_MEM_D_PINLOC_35                               = 0,
   parameter PORT_MEM_D_PINLOC_36                               = 0,
   parameter PORT_MEM_D_PINLOC_37                               = 0,
   parameter PORT_MEM_D_PINLOC_38                               = 0,
   parameter PORT_MEM_D_PINLOC_39                               = 0,
   parameter PORT_MEM_D_PINLOC_40                               = 0,
   parameter PORT_MEM_D_PINLOC_41                               = 0,
   parameter PORT_MEM_D_PINLOC_42                               = 0,
   parameter PORT_MEM_D_PINLOC_43                               = 0,
   parameter PORT_MEM_D_PINLOC_44                               = 0,
   parameter PORT_MEM_D_PINLOC_45                               = 0,
   parameter PORT_MEM_D_PINLOC_46                               = 0,
   parameter PORT_MEM_D_PINLOC_47                               = 0,
   parameter PORT_MEM_D_PINLOC_48                               = 0,
   parameter PORT_MEM_D_PINLOC_AUTOGEN_WCNT                     = 0,
   parameter PORT_MEM_DQ_WIDTH                                  = 0,
   parameter PORT_MEM_DQ_PINLOC_0                               = 0,
   parameter PORT_MEM_DQ_PINLOC_1                               = 0,
   parameter PORT_MEM_DQ_PINLOC_2                               = 0,
   parameter PORT_MEM_DQ_PINLOC_3                               = 0,
   parameter PORT_MEM_DQ_PINLOC_4                               = 0,
   parameter PORT_MEM_DQ_PINLOC_5                               = 0,
   parameter PORT_MEM_DQ_PINLOC_6                               = 0,
   parameter PORT_MEM_DQ_PINLOC_7                               = 0,
   parameter PORT_MEM_DQ_PINLOC_8                               = 0,
   parameter PORT_MEM_DQ_PINLOC_9                               = 0,
   parameter PORT_MEM_DQ_PINLOC_10                              = 0,
   parameter PORT_MEM_DQ_PINLOC_11                              = 0,
   parameter PORT_MEM_DQ_PINLOC_12                              = 0,
   parameter PORT_MEM_DQ_PINLOC_13                              = 0,
   parameter PORT_MEM_DQ_PINLOC_14                              = 0,
   parameter PORT_MEM_DQ_PINLOC_15                              = 0,
   parameter PORT_MEM_DQ_PINLOC_16                              = 0,
   parameter PORT_MEM_DQ_PINLOC_17                              = 0,
   parameter PORT_MEM_DQ_PINLOC_18                              = 0,
   parameter PORT_MEM_DQ_PINLOC_19                              = 0,
   parameter PORT_MEM_DQ_PINLOC_20                              = 0,
   parameter PORT_MEM_DQ_PINLOC_21                              = 0,
   parameter PORT_MEM_DQ_PINLOC_22                              = 0,
   parameter PORT_MEM_DQ_PINLOC_23                              = 0,
   parameter PORT_MEM_DQ_PINLOC_24                              = 0,
   parameter PORT_MEM_DQ_PINLOC_25                              = 0,
   parameter PORT_MEM_DQ_PINLOC_26                              = 0,
   parameter PORT_MEM_DQ_PINLOC_27                              = 0,
   parameter PORT_MEM_DQ_PINLOC_28                              = 0,
   parameter PORT_MEM_DQ_PINLOC_29                              = 0,
   parameter PORT_MEM_DQ_PINLOC_30                              = 0,
   parameter PORT_MEM_DQ_PINLOC_31                              = 0,
   parameter PORT_MEM_DQ_PINLOC_32                              = 0,
   parameter PORT_MEM_DQ_PINLOC_33                              = 0,
   parameter PORT_MEM_DQ_PINLOC_34                              = 0,
   parameter PORT_MEM_DQ_PINLOC_35                              = 0,
   parameter PORT_MEM_DQ_PINLOC_36                              = 0,
   parameter PORT_MEM_DQ_PINLOC_37                              = 0,
   parameter PORT_MEM_DQ_PINLOC_38                              = 0,
   parameter PORT_MEM_DQ_PINLOC_39                              = 0,
   parameter PORT_MEM_DQ_PINLOC_40                              = 0,
   parameter PORT_MEM_DQ_PINLOC_41                              = 0,
   parameter PORT_MEM_DQ_PINLOC_42                              = 0,
   parameter PORT_MEM_DQ_PINLOC_43                              = 0,
   parameter PORT_MEM_DQ_PINLOC_44                              = 0,
   parameter PORT_MEM_DQ_PINLOC_45                              = 0,
   parameter PORT_MEM_DQ_PINLOC_46                              = 0,
   parameter PORT_MEM_DQ_PINLOC_47                              = 0,
   parameter PORT_MEM_DQ_PINLOC_48                              = 0,
   parameter PORT_MEM_DQ_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_DBI_N_WIDTH                               = 0,
   parameter PORT_MEM_DBI_N_PINLOC_0                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_1                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_2                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_3                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_4                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_5                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_6                            = 0,
   parameter PORT_MEM_DBI_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_DQA_WIDTH                                 = 0,
   parameter PORT_MEM_DQA_PINLOC_0                              = 0,
   parameter PORT_MEM_DQA_PINLOC_1                              = 0,
   parameter PORT_MEM_DQA_PINLOC_2                              = 0,
   parameter PORT_MEM_DQA_PINLOC_3                              = 0,
   parameter PORT_MEM_DQA_PINLOC_4                              = 0,
   parameter PORT_MEM_DQA_PINLOC_5                              = 0,
   parameter PORT_MEM_DQA_PINLOC_6                              = 0,
   parameter PORT_MEM_DQA_PINLOC_7                              = 0,
   parameter PORT_MEM_DQA_PINLOC_8                              = 0,
   parameter PORT_MEM_DQA_PINLOC_9                              = 0,
   parameter PORT_MEM_DQA_PINLOC_10                             = 0,
   parameter PORT_MEM_DQA_PINLOC_11                             = 0,
   parameter PORT_MEM_DQA_PINLOC_12                             = 0,
   parameter PORT_MEM_DQA_PINLOC_13                             = 0,
   parameter PORT_MEM_DQA_PINLOC_14                             = 0,
   parameter PORT_MEM_DQA_PINLOC_15                             = 0,
   parameter PORT_MEM_DQA_PINLOC_16                             = 0,
   parameter PORT_MEM_DQA_PINLOC_17                             = 0,
   parameter PORT_MEM_DQA_PINLOC_18                             = 0,
   parameter PORT_MEM_DQA_PINLOC_19                             = 0,
   parameter PORT_MEM_DQA_PINLOC_20                             = 0,
   parameter PORT_MEM_DQA_PINLOC_21                             = 0,
   parameter PORT_MEM_DQA_PINLOC_22                             = 0,
   parameter PORT_MEM_DQA_PINLOC_23                             = 0,
   parameter PORT_MEM_DQA_PINLOC_24                             = 0,
   parameter PORT_MEM_DQA_PINLOC_25                             = 0,
   parameter PORT_MEM_DQA_PINLOC_26                             = 0,
   parameter PORT_MEM_DQA_PINLOC_27                             = 0,
   parameter PORT_MEM_DQA_PINLOC_28                             = 0,
   parameter PORT_MEM_DQA_PINLOC_29                             = 0,
   parameter PORT_MEM_DQA_PINLOC_30                             = 0,
   parameter PORT_MEM_DQA_PINLOC_31                             = 0,
   parameter PORT_MEM_DQA_PINLOC_32                             = 0,
   parameter PORT_MEM_DQA_PINLOC_33                             = 0,
   parameter PORT_MEM_DQA_PINLOC_34                             = 0,
   parameter PORT_MEM_DQA_PINLOC_35                             = 0,
   parameter PORT_MEM_DQA_PINLOC_36                             = 0,
   parameter PORT_MEM_DQA_PINLOC_37                             = 0,
   parameter PORT_MEM_DQA_PINLOC_38                             = 0,
   parameter PORT_MEM_DQA_PINLOC_39                             = 0,
   parameter PORT_MEM_DQA_PINLOC_40                             = 0,
   parameter PORT_MEM_DQA_PINLOC_41                             = 0,
   parameter PORT_MEM_DQA_PINLOC_42                             = 0,
   parameter PORT_MEM_DQA_PINLOC_43                             = 0,
   parameter PORT_MEM_DQA_PINLOC_44                             = 0,
   parameter PORT_MEM_DQA_PINLOC_45                             = 0,
   parameter PORT_MEM_DQA_PINLOC_46                             = 0,
   parameter PORT_MEM_DQA_PINLOC_47                             = 0,
   parameter PORT_MEM_DQA_PINLOC_48                             = 0,
   parameter PORT_MEM_DQA_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_DQB_WIDTH                                 = 0,
   parameter PORT_MEM_DQB_PINLOC_0                              = 0,
   parameter PORT_MEM_DQB_PINLOC_1                              = 0,
   parameter PORT_MEM_DQB_PINLOC_2                              = 0,
   parameter PORT_MEM_DQB_PINLOC_3                              = 0,
   parameter PORT_MEM_DQB_PINLOC_4                              = 0,
   parameter PORT_MEM_DQB_PINLOC_5                              = 0,
   parameter PORT_MEM_DQB_PINLOC_6                              = 0,
   parameter PORT_MEM_DQB_PINLOC_7                              = 0,
   parameter PORT_MEM_DQB_PINLOC_8                              = 0,
   parameter PORT_MEM_DQB_PINLOC_9                              = 0,
   parameter PORT_MEM_DQB_PINLOC_10                             = 0,
   parameter PORT_MEM_DQB_PINLOC_11                             = 0,
   parameter PORT_MEM_DQB_PINLOC_12                             = 0,
   parameter PORT_MEM_DQB_PINLOC_13                             = 0,
   parameter PORT_MEM_DQB_PINLOC_14                             = 0,
   parameter PORT_MEM_DQB_PINLOC_15                             = 0,
   parameter PORT_MEM_DQB_PINLOC_16                             = 0,
   parameter PORT_MEM_DQB_PINLOC_17                             = 0,
   parameter PORT_MEM_DQB_PINLOC_18                             = 0,
   parameter PORT_MEM_DQB_PINLOC_19                             = 0,
   parameter PORT_MEM_DQB_PINLOC_20                             = 0,
   parameter PORT_MEM_DQB_PINLOC_21                             = 0,
   parameter PORT_MEM_DQB_PINLOC_22                             = 0,
   parameter PORT_MEM_DQB_PINLOC_23                             = 0,
   parameter PORT_MEM_DQB_PINLOC_24                             = 0,
   parameter PORT_MEM_DQB_PINLOC_25                             = 0,
   parameter PORT_MEM_DQB_PINLOC_26                             = 0,
   parameter PORT_MEM_DQB_PINLOC_27                             = 0,
   parameter PORT_MEM_DQB_PINLOC_28                             = 0,
   parameter PORT_MEM_DQB_PINLOC_29                             = 0,
   parameter PORT_MEM_DQB_PINLOC_30                             = 0,
   parameter PORT_MEM_DQB_PINLOC_31                             = 0,
   parameter PORT_MEM_DQB_PINLOC_32                             = 0,
   parameter PORT_MEM_DQB_PINLOC_33                             = 0,
   parameter PORT_MEM_DQB_PINLOC_34                             = 0,
   parameter PORT_MEM_DQB_PINLOC_35                             = 0,
   parameter PORT_MEM_DQB_PINLOC_36                             = 0,
   parameter PORT_MEM_DQB_PINLOC_37                             = 0,
   parameter PORT_MEM_DQB_PINLOC_38                             = 0,
   parameter PORT_MEM_DQB_PINLOC_39                             = 0,
   parameter PORT_MEM_DQB_PINLOC_40                             = 0,
   parameter PORT_MEM_DQB_PINLOC_41                             = 0,
   parameter PORT_MEM_DQB_PINLOC_42                             = 0,
   parameter PORT_MEM_DQB_PINLOC_43                             = 0,
   parameter PORT_MEM_DQB_PINLOC_44                             = 0,
   parameter PORT_MEM_DQB_PINLOC_45                             = 0,
   parameter PORT_MEM_DQB_PINLOC_46                             = 0,
   parameter PORT_MEM_DQB_PINLOC_47                             = 0,
   parameter PORT_MEM_DQB_PINLOC_48                             = 0,
   parameter PORT_MEM_DQB_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_DINVA_WIDTH                               = 0,
   parameter PORT_MEM_DINVA_PINLOC_0                            = 0,
   parameter PORT_MEM_DINVA_PINLOC_1                            = 0,
   parameter PORT_MEM_DINVA_PINLOC_2                            = 0,
   parameter PORT_MEM_DINVA_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_DINVB_WIDTH                               = 0,
   parameter PORT_MEM_DINVB_PINLOC_0                            = 0,
   parameter PORT_MEM_DINVB_PINLOC_1                            = 0,
   parameter PORT_MEM_DINVB_PINLOC_2                            = 0,
   parameter PORT_MEM_DINVB_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_Q_WIDTH                                   = 0,
   parameter PORT_MEM_Q_PINLOC_0                                = 0,
   parameter PORT_MEM_Q_PINLOC_1                                = 0,
   parameter PORT_MEM_Q_PINLOC_2                                = 0,
   parameter PORT_MEM_Q_PINLOC_3                                = 0,
   parameter PORT_MEM_Q_PINLOC_4                                = 0,
   parameter PORT_MEM_Q_PINLOC_5                                = 0,
   parameter PORT_MEM_Q_PINLOC_6                                = 0,
   parameter PORT_MEM_Q_PINLOC_7                                = 0,
   parameter PORT_MEM_Q_PINLOC_8                                = 0,
   parameter PORT_MEM_Q_PINLOC_9                                = 0,
   parameter PORT_MEM_Q_PINLOC_10                               = 0,
   parameter PORT_MEM_Q_PINLOC_11                               = 0,
   parameter PORT_MEM_Q_PINLOC_12                               = 0,
   parameter PORT_MEM_Q_PINLOC_13                               = 0,
   parameter PORT_MEM_Q_PINLOC_14                               = 0,
   parameter PORT_MEM_Q_PINLOC_15                               = 0,
   parameter PORT_MEM_Q_PINLOC_16                               = 0,
   parameter PORT_MEM_Q_PINLOC_17                               = 0,
   parameter PORT_MEM_Q_PINLOC_18                               = 0,
   parameter PORT_MEM_Q_PINLOC_19                               = 0,
   parameter PORT_MEM_Q_PINLOC_20                               = 0,
   parameter PORT_MEM_Q_PINLOC_21                               = 0,
   parameter PORT_MEM_Q_PINLOC_22                               = 0,
   parameter PORT_MEM_Q_PINLOC_23                               = 0,
   parameter PORT_MEM_Q_PINLOC_24                               = 0,
   parameter PORT_MEM_Q_PINLOC_25                               = 0,
   parameter PORT_MEM_Q_PINLOC_26                               = 0,
   parameter PORT_MEM_Q_PINLOC_27                               = 0,
   parameter PORT_MEM_Q_PINLOC_28                               = 0,
   parameter PORT_MEM_Q_PINLOC_29                               = 0,
   parameter PORT_MEM_Q_PINLOC_30                               = 0,
   parameter PORT_MEM_Q_PINLOC_31                               = 0,
   parameter PORT_MEM_Q_PINLOC_32                               = 0,
   parameter PORT_MEM_Q_PINLOC_33                               = 0,
   parameter PORT_MEM_Q_PINLOC_34                               = 0,
   parameter PORT_MEM_Q_PINLOC_35                               = 0,
   parameter PORT_MEM_Q_PINLOC_36                               = 0,
   parameter PORT_MEM_Q_PINLOC_37                               = 0,
   parameter PORT_MEM_Q_PINLOC_38                               = 0,
   parameter PORT_MEM_Q_PINLOC_39                               = 0,
   parameter PORT_MEM_Q_PINLOC_40                               = 0,
   parameter PORT_MEM_Q_PINLOC_41                               = 0,
   parameter PORT_MEM_Q_PINLOC_42                               = 0,
   parameter PORT_MEM_Q_PINLOC_43                               = 0,
   parameter PORT_MEM_Q_PINLOC_44                               = 0,
   parameter PORT_MEM_Q_PINLOC_45                               = 0,
   parameter PORT_MEM_Q_PINLOC_46                               = 0,
   parameter PORT_MEM_Q_PINLOC_47                               = 0,
   parameter PORT_MEM_Q_PINLOC_48                               = 0,
   parameter PORT_MEM_Q_PINLOC_AUTOGEN_WCNT                     = 0,
   parameter PORT_MEM_DQS_WIDTH                                 = 0,
   parameter PORT_MEM_DQS_PINLOC_0                              = 0,
   parameter PORT_MEM_DQS_PINLOC_1                              = 0,
   parameter PORT_MEM_DQS_PINLOC_2                              = 0,
   parameter PORT_MEM_DQS_PINLOC_3                              = 0,
   parameter PORT_MEM_DQS_PINLOC_4                              = 0,
   parameter PORT_MEM_DQS_PINLOC_5                              = 0,
   parameter PORT_MEM_DQS_PINLOC_6                              = 0,
   parameter PORT_MEM_DQS_PINLOC_7                              = 0,
   parameter PORT_MEM_DQS_PINLOC_8                              = 0,
   parameter PORT_MEM_DQS_PINLOC_9                              = 0,
   parameter PORT_MEM_DQS_PINLOC_10                             = 0,
   parameter PORT_MEM_DQS_PINLOC_11                             = 0,
   parameter PORT_MEM_DQS_PINLOC_12                             = 0,
   parameter PORT_MEM_DQS_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_DQS_N_WIDTH                               = 0,
   parameter PORT_MEM_DQS_N_PINLOC_0                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_1                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_2                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_3                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_4                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_5                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_6                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_7                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_8                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_9                            = 0,
   parameter PORT_MEM_DQS_N_PINLOC_10                           = 0,
   parameter PORT_MEM_DQS_N_PINLOC_11                           = 0,
   parameter PORT_MEM_DQS_N_PINLOC_12                           = 0,
   parameter PORT_MEM_DQS_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_QK_WIDTH                                  = 0,
   parameter PORT_MEM_QK_PINLOC_0                               = 0,
   parameter PORT_MEM_QK_PINLOC_1                               = 0,
   parameter PORT_MEM_QK_PINLOC_2                               = 0,
   parameter PORT_MEM_QK_PINLOC_3                               = 0,
   parameter PORT_MEM_QK_PINLOC_4                               = 0,
   parameter PORT_MEM_QK_PINLOC_5                               = 0,
   parameter PORT_MEM_QK_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_QK_N_WIDTH                                = 0,
   parameter PORT_MEM_QK_N_PINLOC_0                             = 0,
   parameter PORT_MEM_QK_N_PINLOC_1                             = 0,
   parameter PORT_MEM_QK_N_PINLOC_2                             = 0,
   parameter PORT_MEM_QK_N_PINLOC_3                             = 0,
   parameter PORT_MEM_QK_N_PINLOC_4                             = 0,
   parameter PORT_MEM_QK_N_PINLOC_5                             = 0,
   parameter PORT_MEM_QK_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_QKA_WIDTH                                 = 0,
   parameter PORT_MEM_QKA_PINLOC_0                              = 0,
   parameter PORT_MEM_QKA_PINLOC_1                              = 0,
   parameter PORT_MEM_QKA_PINLOC_2                              = 0,
   parameter PORT_MEM_QKA_PINLOC_3                              = 0,
   parameter PORT_MEM_QKA_PINLOC_4                              = 0,
   parameter PORT_MEM_QKA_PINLOC_5                              = 0,
   parameter PORT_MEM_QKA_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_QKA_N_WIDTH                               = 0,
   parameter PORT_MEM_QKA_N_PINLOC_0                            = 0,
   parameter PORT_MEM_QKA_N_PINLOC_1                            = 0,
   parameter PORT_MEM_QKA_N_PINLOC_2                            = 0,
   parameter PORT_MEM_QKA_N_PINLOC_3                            = 0,
   parameter PORT_MEM_QKA_N_PINLOC_4                            = 0,
   parameter PORT_MEM_QKA_N_PINLOC_5                            = 0,
   parameter PORT_MEM_QKA_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_QKB_WIDTH                                 = 0,
   parameter PORT_MEM_QKB_PINLOC_0                              = 0,
   parameter PORT_MEM_QKB_PINLOC_1                              = 0,
   parameter PORT_MEM_QKB_PINLOC_2                              = 0,
   parameter PORT_MEM_QKB_PINLOC_3                              = 0,
   parameter PORT_MEM_QKB_PINLOC_4                              = 0,
   parameter PORT_MEM_QKB_PINLOC_5                              = 0,
   parameter PORT_MEM_QKB_PINLOC_AUTOGEN_WCNT                   = 0,
   parameter PORT_MEM_QKB_N_WIDTH                               = 0,
   parameter PORT_MEM_QKB_N_PINLOC_0                            = 0,
   parameter PORT_MEM_QKB_N_PINLOC_1                            = 0,
   parameter PORT_MEM_QKB_N_PINLOC_2                            = 0,
   parameter PORT_MEM_QKB_N_PINLOC_3                            = 0,
   parameter PORT_MEM_QKB_N_PINLOC_4                            = 0,
   parameter PORT_MEM_QKB_N_PINLOC_5                            = 0,
   parameter PORT_MEM_QKB_N_PINLOC_AUTOGEN_WCNT                 = 0,
   parameter PORT_MEM_CQ_WIDTH                                  = 0,
   parameter PORT_MEM_CQ_PINLOC_0                               = 0,
   parameter PORT_MEM_CQ_PINLOC_1                               = 0,
   parameter PORT_MEM_CQ_PINLOC_AUTOGEN_WCNT                    = 0,
   parameter PORT_MEM_CQ_N_WIDTH                                = 0,
   parameter PORT_MEM_CQ_N_PINLOC_0                             = 0,
   parameter PORT_MEM_CQ_N_PINLOC_1                             = 0,
   parameter PORT_MEM_CQ_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_MEM_ALERT_N_WIDTH                             = 0,
   parameter PORT_MEM_ALERT_N_PINLOC_0                          = 0,
   parameter PORT_MEM_ALERT_N_PINLOC_1                          = 0,
   parameter PORT_MEM_ALERT_N_PINLOC_AUTOGEN_WCNT               = 0,
   parameter PORT_MEM_PE_N_WIDTH                                = 0,
   parameter PORT_MEM_PE_N_PINLOC_0                             = 0,
   parameter PORT_MEM_PE_N_PINLOC_1                             = 0,
   parameter PORT_MEM_PE_N_PINLOC_AUTOGEN_WCNT                  = 0,
   parameter PORT_CLKS_SHARING_MASTER_OUT_WIDTH                 = 0,
   parameter PORT_CLKS_SHARING_SLAVE_IN_WIDTH                   = 0,
   parameter PORT_AFI_RLAT_WIDTH                                = 0,
   parameter PORT_AFI_WLAT_WIDTH                                = 0,
   parameter PORT_AFI_SEQ_BUSY_WIDTH                            = 0,
   parameter PORT_AFI_ADDR_WIDTH                                = 0,
   parameter PORT_AFI_BA_WIDTH                                  = 0,
   parameter PORT_AFI_BG_WIDTH                                  = 0,
   parameter PORT_AFI_C_WIDTH                                   = 0,
   parameter PORT_AFI_CKE_WIDTH                                 = 0,
   parameter PORT_AFI_CS_N_WIDTH                                = 0,
   parameter PORT_AFI_RM_WIDTH                                  = 0,
   parameter PORT_AFI_ODT_WIDTH                                 = 0,
   parameter PORT_AFI_RAS_N_WIDTH                               = 0,
   parameter PORT_AFI_CAS_N_WIDTH                               = 0,
   parameter PORT_AFI_WE_N_WIDTH                                = 0,
   parameter PORT_AFI_RST_N_WIDTH                               = 0,
   parameter PORT_AFI_ACT_N_WIDTH                               = 0,
   parameter PORT_AFI_PAR_WIDTH                                 = 0,
   parameter PORT_AFI_CA_WIDTH                                  = 0,
   parameter PORT_AFI_REF_N_WIDTH                               = 0,
   parameter PORT_AFI_WPS_N_WIDTH                               = 0,
   parameter PORT_AFI_RPS_N_WIDTH                               = 0,
   parameter PORT_AFI_DOFF_N_WIDTH                              = 0,
   parameter PORT_AFI_LD_N_WIDTH                                = 0,
   parameter PORT_AFI_RW_N_WIDTH                                = 0,
   parameter PORT_AFI_LBK0_N_WIDTH                              = 0,
   parameter PORT_AFI_LBK1_N_WIDTH                              = 0,
   parameter PORT_AFI_CFG_N_WIDTH                               = 0,
   parameter PORT_AFI_AP_WIDTH                                  = 0,
   parameter PORT_AFI_AINV_WIDTH                                = 0,
   parameter PORT_AFI_DM_WIDTH                                  = 0,
   parameter PORT_AFI_DM_N_WIDTH                                = 0,
   parameter PORT_AFI_BWS_N_WIDTH                               = 0,
   parameter PORT_AFI_RDATA_DBI_N_WIDTH                         = 0,
   parameter PORT_AFI_WDATA_DBI_N_WIDTH                         = 0,
   parameter PORT_AFI_RDATA_DINV_WIDTH                          = 0,
   parameter PORT_AFI_WDATA_DINV_WIDTH                          = 0,
   parameter PORT_AFI_DQS_BURST_WIDTH                           = 0,
   parameter PORT_AFI_WDATA_VALID_WIDTH                         = 0,
   parameter PORT_AFI_WDATA_WIDTH                               = 0,
   parameter PORT_AFI_RDATA_EN_FULL_WIDTH                       = 0,
   parameter PORT_AFI_RDATA_WIDTH                               = 0,
   parameter PORT_AFI_RDATA_VALID_WIDTH                         = 0,
   parameter PORT_AFI_RRANK_WIDTH                               = 0,
   parameter PORT_AFI_WRANK_WIDTH                               = 0,
   parameter PORT_AFI_ALERT_N_WIDTH                             = 0,
   parameter PORT_AFI_PE_N_WIDTH                                = 0,
   parameter PORT_CTRL_AST_CMD_DATA_WIDTH                       = 0,
   parameter PORT_CTRL_AST_WR_DATA_WIDTH                        = 0,
   parameter PORT_CTRL_AST_RD_DATA_WIDTH                        = 0,
   parameter PORT_CTRL_AMM_ADDRESS_WIDTH                        = 0,
   parameter PORT_CTRL_AMM_RDATA_WIDTH                          = 0,
   parameter PORT_CTRL_AMM_WDATA_WIDTH                          = 0,
   parameter PORT_CTRL_AMM_BCOUNT_WIDTH                         = 0,
   parameter PORT_CTRL_AMM_BYTEEN_WIDTH                         = 0,
   parameter PORT_CTRL_USER_REFRESH_REQ_WIDTH                   = 0,
   parameter PORT_CTRL_USER_REFRESH_BANK_WIDTH                  = 0,
   parameter PORT_CTRL_SELF_REFRESH_REQ_WIDTH                   = 0,
   parameter PORT_CTRL_ECC_WRITE_INFO_WIDTH                     = 0,
   parameter PORT_CTRL_ECC_RDATA_ID_WIDTH                       = 0,
   parameter PORT_CTRL_ECC_READ_INFO_WIDTH                      = 0,
   parameter PORT_CTRL_ECC_CMD_INFO_WIDTH                       = 0,
   parameter PORT_CTRL_ECC_WB_POINTER_WIDTH                     = 0,
   parameter PORT_CTRL_MMR_SLAVE_ADDRESS_WIDTH                  = 0,
   parameter PORT_CTRL_MMR_SLAVE_RDATA_WIDTH                    = 0,
   parameter PORT_CTRL_MMR_SLAVE_WDATA_WIDTH                    = 0,
   parameter PORT_CTRL_MMR_SLAVE_BCOUNT_WIDTH                   = 0,
   parameter PORT_HPS_EMIF_H2E_WIDTH                            = 0,
   parameter PORT_HPS_EMIF_E2H_WIDTH                            = 0,
   parameter PORT_HPS_EMIF_H2E_GP_WIDTH                         = 0,
   parameter PORT_HPS_EMIF_E2H_GP_WIDTH                         = 0,
   parameter PORT_CAL_DEBUG_ADDRESS_WIDTH                       = 0,
   parameter PORT_CAL_DEBUG_RDATA_WIDTH                         = 0,
   parameter PORT_CAL_DEBUG_WDATA_WIDTH                         = 0,
   parameter PORT_CAL_DEBUG_BYTEEN_WIDTH                        = 0,
   parameter PORT_CAL_DEBUG_OUT_ADDRESS_WIDTH                   = 0,
   parameter PORT_CAL_DEBUG_OUT_RDATA_WIDTH                     = 0,
   parameter PORT_CAL_DEBUG_OUT_WDATA_WIDTH                     = 0,
   parameter PORT_CAL_DEBUG_OUT_BYTEEN_WIDTH                    = 0,
   parameter PORT_CAL_MASTER_ADDRESS_WIDTH                      = 0,
   parameter PORT_CAL_MASTER_RDATA_WIDTH                        = 0,
   parameter PORT_CAL_MASTER_WDATA_WIDTH                        = 0,
   parameter PORT_CAL_MASTER_BYTEEN_WIDTH                       = 0,
   parameter PORT_DFT_NF_IOAUX_PIO_IN_WIDTH                     = 0,
   parameter PORT_DFT_NF_IOAUX_PIO_OUT_WIDTH                    = 0,
   parameter PORT_DFT_NF_PA_DPRIO_REG_ADDR_WIDTH                = 0,
   parameter PORT_DFT_NF_PA_DPRIO_WRITEDATA_WIDTH               = 0,
   parameter PORT_DFT_NF_PA_DPRIO_READDATA_WIDTH                = 0,
   parameter PORT_DFT_NF_PLL_CNTSEL_WIDTH                       = 0,
   parameter PORT_DFT_NF_PLL_NUM_SHIFT_WIDTH                    = 0,
   parameter PORT_DFT_NF_CORE_CLK_BUF_OUT_WIDTH                 = 0,
   parameter PORT_DFT_NF_CORE_CLK_LOCKED_WIDTH                  = 0,
   parameter PLL_VCO_FREQ_MHZ_INT                               = 0,
   parameter PLL_VCO_TO_MEM_CLK_FREQ_RATIO                      = 0,
   parameter PLL_PHY_CLK_VCO_PHASE                              = 0,
   parameter PLL_VCO_FREQ_PS_STR                                = "",
   parameter PLL_REF_CLK_FREQ_PS_STR                            = "",
   parameter PLL_REF_CLK_FREQ_PS                                = 0,
   parameter PLL_SIM_VCO_FREQ_PS                                = 0,
   parameter PLL_SIM_PHYCLK_0_FREQ_PS                           = 0,
   parameter PLL_SIM_PHYCLK_1_FREQ_PS                           = 0,
   parameter PLL_SIM_PHYCLK_FB_FREQ_PS                          = 0,
   parameter PLL_SIM_PHY_CLK_VCO_PHASE_PS                       = 0,
   parameter PLL_SIM_CAL_SLAVE_CLK_FREQ_PS                      = 0,
   parameter PLL_SIM_CAL_MASTER_CLK_FREQ_PS                     = 0,
   parameter PLL_M_CNT_HIGH                                     = 0,
   parameter PLL_M_CNT_LOW                                      = 0,
   parameter PLL_N_CNT_HIGH                                     = 0,
   parameter PLL_N_CNT_LOW                                      = 0,
   parameter PLL_M_CNT_BYPASS_EN                                = "",
   parameter PLL_N_CNT_BYPASS_EN                                = "",
   parameter PLL_M_CNT_EVEN_DUTY_EN                             = "",
   parameter PLL_N_CNT_EVEN_DUTY_EN                             = "",
   parameter PLL_FBCLK_MUX_1                                    = "",
   parameter PLL_FBCLK_MUX_2                                    = "",
   parameter PLL_M_CNT_IN_SRC                                   = "",
   parameter PLL_CP_SETTING                                     = "",
   parameter PLL_BW_CTRL                                        = "",
   parameter PLL_BW_SEL                                         = "",
   parameter PLL_C_CNT_HIGH_0                                   = 0,
   parameter PLL_C_CNT_LOW_0                                    = 0,
   parameter PLL_C_CNT_PRST_0                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_0                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_0                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_0                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_0                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_0                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_0                             = 0,
   parameter PLL_C_CNT_OUT_EN_0                                 = "",
   parameter PLL_C_CNT_HIGH_1                                   = 0,
   parameter PLL_C_CNT_LOW_1                                    = 0,
   parameter PLL_C_CNT_PRST_1                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_1                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_1                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_1                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_1                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_1                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_1                             = 0,
   parameter PLL_C_CNT_OUT_EN_1                                 = "",
   parameter PLL_C_CNT_HIGH_2                                   = 0,
   parameter PLL_C_CNT_LOW_2                                    = 0,
   parameter PLL_C_CNT_PRST_2                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_2                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_2                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_2                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_2                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_2                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_2                             = 0,
   parameter PLL_C_CNT_OUT_EN_2                                 = "",
   parameter PLL_C_CNT_HIGH_3                                   = 0,
   parameter PLL_C_CNT_LOW_3                                    = 0,
   parameter PLL_C_CNT_PRST_3                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_3                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_3                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_3                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_3                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_3                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_3                             = 0,
   parameter PLL_C_CNT_OUT_EN_3                                 = "",
   parameter PLL_C_CNT_HIGH_4                                   = 0,
   parameter PLL_C_CNT_LOW_4                                    = 0,
   parameter PLL_C_CNT_PRST_4                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_4                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_4                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_4                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_4                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_4                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_4                             = 0,
   parameter PLL_C_CNT_OUT_EN_4                                 = "",
   parameter PLL_C_CNT_HIGH_5                                   = 0,
   parameter PLL_C_CNT_LOW_5                                    = 0,
   parameter PLL_C_CNT_PRST_5                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_5                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_5                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_5                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_5                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_5                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_5                             = 0,
   parameter PLL_C_CNT_OUT_EN_5                                 = "",
   parameter PLL_C_CNT_HIGH_6                                   = 0,
   parameter PLL_C_CNT_LOW_6                                    = 0,
   parameter PLL_C_CNT_PRST_6                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_6                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_6                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_6                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_6                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_6                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_6                             = 0,
   parameter PLL_C_CNT_OUT_EN_6                                 = "",
   parameter PLL_C_CNT_HIGH_7                                   = 0,
   parameter PLL_C_CNT_LOW_7                                    = 0,
   parameter PLL_C_CNT_PRST_7                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_7                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_7                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_7                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_7                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_7                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_7                             = 0,
   parameter PLL_C_CNT_OUT_EN_7                                 = "",
   parameter PLL_C_CNT_HIGH_8                                   = 0,
   parameter PLL_C_CNT_LOW_8                                    = 0,
   parameter PLL_C_CNT_PRST_8                                   = 0,
   parameter PLL_C_CNT_PH_MUX_PRST_8                            = 0,
   parameter PLL_C_CNT_BYPASS_EN_8                              = "",
   parameter PLL_C_CNT_EVEN_DUTY_EN_8                           = "",
   parameter PLL_C_CNT_FREQ_PS_STR_8                            = "",
   parameter PLL_C_CNT_PHASE_PS_STR_8                           = "",
   parameter PLL_C_CNT_DUTY_CYCLE_8                             = 0,
   parameter PLL_C_CNT_OUT_EN_8                                 = ""
) (
   input  logic            global_reset_n,
   input  logic            pll_ref_clk,
   output logic            pll_locked,
   output logic            pll_extra_clk_0,
   output logic            pll_extra_clk_1,
   output logic            pll_extra_clk_2,
   output logic            pll_extra_clk_3,
   input  logic            oct_rzqin,
   output logic [0:0]      mem_ck,
   output logic [0:0]      mem_ck_n,
   output logic [16:0]     mem_a,
   output logic [0:0]      mem_act_n,
   output logic [1:0]      mem_ba,
   output logic [1:0]      mem_bg,
   output logic [0:0]      mem_c,
   output logic [0:0]      mem_cke,
   output logic [0:0]      mem_cs_n,
   output logic [0:0]      mem_rm,
   output logic [0:0]      mem_odt,
   output logic [0:0]      mem_reset_n,
   output logic [0:0]      mem_par,
   input  logic [0:0]      mem_alert_n,
   inout  tri   [7:0]      mem_dqs,
   inout  tri   [7:0]      mem_dqs_n,
   inout  tri   [63:0]     mem_dq,
   inout  tri   [7:0]      mem_dbi_n,
   output logic [0:0]      mem_dk,
   output logic [0:0]      mem_dk_n,
   output logic [0:0]      mem_dka,
   output logic [0:0]      mem_dka_n,
   output logic [0:0]      mem_dkb,
   output logic [0:0]      mem_dkb_n,
   output logic [0:0]      mem_k,
   output logic [0:0]      mem_k_n,
   output logic [0:0]      mem_ras_n,
   output logic [0:0]      mem_cas_n,
   output logic [0:0]      mem_we_n,
   output logic [0:0]      mem_ca,
   output logic [0:0]      mem_ref_n,
   output logic [0:0]      mem_wps_n,
   output logic [0:0]      mem_rps_n,
   output logic [0:0]      mem_doff_n,
   output logic [0:0]      mem_lda_n,
   output logic [0:0]      mem_ldb_n,
   output logic [0:0]      mem_rwa_n,
   output logic [0:0]      mem_rwb_n,
   output logic [0:0]      mem_lbk0_n,
   output logic [0:0]      mem_lbk1_n,
   output logic [0:0]      mem_cfg_n,
   output logic [0:0]      mem_ap,
   output logic [0:0]      mem_ainv,
   output logic [0:0]      mem_dm,
   output logic [0:0]      mem_bws_n,
   output logic [0:0]      mem_d,
   inout  tri   [0:0]      mem_dqa,
   inout  tri   [0:0]      mem_dqb,
   inout  tri   [0:0]      mem_dinva,
   inout  tri   [0:0]      mem_dinvb,
   input  logic [0:0]      mem_q,
   input  logic [0:0]      mem_qk,
   input  logic [0:0]      mem_qk_n,
   input  logic [0:0]      mem_qka,
   input  logic [0:0]      mem_qka_n,
   input  logic [0:0]      mem_qkb,
   input  logic [0:0]      mem_qkb_n,
   input  logic [0:0]      mem_cq,
   input  logic [0:0]      mem_cq_n,
   input  logic [0:0]      mem_pe_n,
   output logic            local_cal_success,
   output logic            local_cal_fail,
   input  logic            vid_cal_done_persist,
   output logic            afi_reset_n,
   output logic            afi_clk,
   output logic            afi_half_clk,
   output logic            emif_usr_reset_n,
   output logic            emif_usr_clk,
   output logic            emif_usr_half_clk,
   output logic            emif_usr_reset_n_sec,
   output logic            emif_usr_clk_sec,
   output logic            emif_usr_half_clk_sec,
   output logic            cal_master_reset_n,
   output logic            cal_master_clk,
   output logic            cal_slave_reset_n,
   output logic            cal_slave_clk,
   input  logic            cal_slave_reset_n_in,
   input  logic            cal_slave_clk_in,
   input  logic            cal_debug_reset_n,
   input  logic            cal_debug_clk,
   output logic            cal_debug_out_reset_n,
   output logic            cal_debug_out_clk,
   output logic [31:0]     clks_sharing_master_out,
   input  logic [31:0]     clks_sharing_slave_in,
   output logic            afi_cal_success,
   output logic            afi_cal_fail,
   input  logic            afi_cal_req,
   output logic [5:0]      afi_rlat,
   output logic [5:0]      afi_wlat,
   output logic [3:0]      afi_seq_busy,
   input  logic            afi_ctl_refresh_done,
   input  logic            afi_ctl_long_idle,
   input  logic            afi_mps_req,
   output logic            afi_mps_ack,
   input  logic [0:0]      afi_addr,
   input  logic [0:0]      afi_ba,
   input  logic [0:0]      afi_bg,
   input  logic [0:0]      afi_c,
   input  logic [0:0]      afi_cke,
   input  logic [0:0]      afi_cs_n,
   input  logic [0:0]      afi_rm,
   input  logic [0:0]      afi_odt,
   input  logic [0:0]      afi_ras_n,
   input  logic [0:0]      afi_cas_n,
   input  logic [0:0]      afi_we_n,
   input  logic [0:0]      afi_rst_n,
   input  logic [0:0]      afi_act_n,
   input  logic [0:0]      afi_par,
   input  logic [0:0]      afi_ca,
   input  logic [0:0]      afi_ref_n,
   input  logic [0:0]      afi_wps_n,
   input  logic [0:0]      afi_rps_n,
   input  logic [0:0]      afi_doff_n,
   input  logic [0:0]      afi_ld_n,
   input  logic [0:0]      afi_rw_n,
   input  logic [0:0]      afi_lbk0_n,
   input  logic [0:0]      afi_lbk1_n,
   input  logic [0:0]      afi_cfg_n,
   input  logic [0:0]      afi_ap,
   input  logic [0:0]      afi_ainv,
   input  logic [0:0]      afi_dm,
   input  logic [0:0]      afi_dm_n,
   input  logic [0:0]      afi_bws_n,
   output logic [0:0]      afi_rdata_dbi_n,
   input  logic [0:0]      afi_wdata_dbi_n,
   output logic [0:0]      afi_rdata_dinv,
   input  logic [0:0]      afi_wdata_dinv,
   input  logic [0:0]      afi_dqs_burst,
   input  logic [0:0]      afi_wdata_valid,
   input  logic [0:0]      afi_wdata,
   input  logic [0:0]      afi_rdata_en_full,
   output logic [0:0]      afi_rdata,
   output logic [0:0]      afi_rdata_valid,
   input  logic [0:0]      afi_rrank,
   input  logic [0:0]      afi_wrank,
   output logic [0:0]      afi_alert_n,
   output logic [0:0]      afi_pe_n,
   input  logic [0:0]      ast_cmd_data_0,
   input  logic            ast_cmd_valid_0,
   output logic            ast_cmd_ready_0,
   input  logic [0:0]      ast_cmd_data_1,
   input  logic            ast_cmd_valid_1,
   output logic            ast_cmd_ready_1,
   input  logic [0:0]      ast_wr_data_0,
   input  logic            ast_wr_valid_0,
   output logic            ast_wr_ready_0,
   input  logic [0:0]      ast_wr_data_1,
   input  logic            ast_wr_valid_1,
   output logic            ast_wr_ready_1,
   output logic [0:0]      ast_rd_data_0,
   output logic            ast_rd_valid_0,
   input  logic            ast_rd_ready_0,
   output logic [0:0]      ast_rd_data_1,
   output logic            ast_rd_valid_1,
   input  logic            ast_rd_ready_1,
   output logic            amm_ready_0,
   input  logic            amm_read_0,
   input  logic            amm_write_0,
   input  logic [25:0]     amm_address_0,
   output logic [511:0]    amm_readdata_0,
   input  logic [511:0]    amm_writedata_0,
   input  logic [6:0]      amm_burstcount_0,
   input  logic [63:0]     amm_byteenable_0,
   input  logic            amm_beginbursttransfer_0,
   output logic            amm_readdatavalid_0,
   output logic            amm_ready_1,
   input  logic            amm_read_1,
   input  logic            amm_write_1,
   input  logic [25:0]     amm_address_1,
   output logic [511:0]    amm_readdata_1,
   input  logic [511:0]    amm_writedata_1,
   input  logic [6:0]      amm_burstcount_1,
   input  logic [63:0]     amm_byteenable_1,
   input  logic            amm_beginbursttransfer_1,
   output logic            amm_readdatavalid_1,
   input  logic            ctrl_user_priority_hi_0,
   input  logic            ctrl_user_priority_hi_1,
   input  logic            ctrl_auto_precharge_req_0,
   input  logic            ctrl_auto_precharge_req_1,
   input  logic [3:0]      ctrl_user_refresh_req,
   input  logic [15:0]     ctrl_user_refresh_bank,
   output logic            ctrl_user_refresh_ack,
   input  logic [3:0]      ctrl_self_refresh_req,
   output logic            ctrl_self_refresh_ack,
   output logic            ctrl_will_refresh,
   input  logic            ctrl_deep_power_down_req,
   output logic            ctrl_deep_power_down_ack,
   output logic            ctrl_power_down_ack,
   input  logic            ctrl_zq_cal_long_req,
   input  logic            ctrl_zq_cal_short_req,
   output logic            ctrl_zq_cal_ack,
   input  logic [14:0]     ctrl_ecc_write_info_0,
   output logic [12:0]     ctrl_ecc_rdata_id_0,
   output logic [2:0]      ctrl_ecc_read_info_0,
   output logic [2:0]      ctrl_ecc_cmd_info_0,
   output logic            ctrl_ecc_idle_0,
   output logic [11:0]     ctrl_ecc_wr_pointer_info_0,
   input  logic [14:0]     ctrl_ecc_write_info_1,
   output logic [12:0]     ctrl_ecc_rdata_id_1,
   output logic [2:0]      ctrl_ecc_read_info_1,
   output logic [2:0]      ctrl_ecc_cmd_info_1,
   output logic            ctrl_ecc_idle_1,
   output logic [11:0]     ctrl_ecc_wr_pointer_info_1,
   output logic            mmr_slave_waitrequest_0,
   input  logic            mmr_slave_read_0,
   input  logic            mmr_slave_write_0,
   input  logic [9:0]      mmr_slave_address_0,
   output logic [31:0]     mmr_slave_readdata_0,
   input  logic [31:0]     mmr_slave_writedata_0,
   input  logic [1:0]      mmr_slave_burstcount_0,
   input  logic            mmr_slave_beginbursttransfer_0,
   output logic            mmr_slave_readdatavalid_0,
   output logic            mmr_slave_waitrequest_1,
   input  logic            mmr_slave_read_1,
   input  logic            mmr_slave_write_1,
   input  logic [9:0]      mmr_slave_address_1,
   output logic [31:0]     mmr_slave_readdata_1,
   input  logic [31:0]     mmr_slave_writedata_1,
   input  logic [1:0]      mmr_slave_burstcount_1,
   input  logic            mmr_slave_beginbursttransfer_1,
   output logic            mmr_slave_readdatavalid_1,
   input  logic [4095:0]   hps_to_emif,
   output logic [4095:0]   emif_to_hps,
   input  logic [1:0]      hps_to_emif_gp,
   output logic [0:0]      emif_to_hps_gp,
   output logic            cal_debug_waitrequest,
   input  logic            cal_debug_read,
   input  logic            cal_debug_write,
   input  logic [23:0]     cal_debug_addr,
   output logic [31:0]     cal_debug_read_data,
   input  logic [31:0]     cal_debug_write_data,
   input  logic [3:0]      cal_debug_byteenable,
   output logic            cal_debug_read_data_valid,
   input  logic            cal_debug_out_waitrequest,
   output logic            cal_debug_out_read,
   output logic            cal_debug_out_write,
   output logic [23:0]     cal_debug_out_addr,
   input  logic [31:0]     cal_debug_out_read_data,
   output logic [31:0]     cal_debug_out_write_data,
   output logic [3:0]      cal_debug_out_byteenable,
   input  logic            cal_debug_out_read_data_valid,
   input  logic            cal_master_waitrequest,
   output logic            cal_master_read,
   output logic            cal_master_write,
   output logic [15:0]     cal_master_addr,
   input  logic [31:0]     cal_master_read_data,
   output logic [31:0]     cal_master_write_data,
   output logic [3:0]      cal_master_byteenable,
   input  logic            cal_master_read_data_valid,
   output logic            cal_master_burstcount,
   output logic            cal_master_debugaccess,
   input  logic [7:0]      ioaux_pio_in,
   output logic [7:0]      ioaux_pio_out,
   input  logic            pa_dprio_clk,
   input  logic            pa_dprio_read,
   input  logic [8:0]      pa_dprio_reg_addr,
   input  logic            pa_dprio_rst_n,
   input  logic            pa_dprio_write,
   input  logic [7:0]      pa_dprio_writedata,
   output logic            pa_dprio_block_select,
   output logic [7:0]      pa_dprio_readdata,
   input  logic            pll_phase_en,
   input  logic            pll_up_dn,
   input  logic [3:0]      pll_cnt_sel,
   input  logic [2:0]      pll_num_phase_shifts,
   output logic            pll_phase_done,
   output logic [1:0]      dft_core_clk_buf_out,
   output logic [1:0]      dft_core_clk_locked
);
   timeunit 1ns;
   timeprecision 1ps;

   emif_ddr4_ddr4b_altera_emif_arch_nf_170_3eabgiq_top # (
      .PROTOCOL_ENUM (PROTOCOL_ENUM),
      .PHY_TARGET_IS_ES (PHY_TARGET_IS_ES),
      .PHY_TARGET_IS_ES2 (PHY_TARGET_IS_ES2),
      .PHY_TARGET_IS_PRODUCTION (PHY_TARGET_IS_PRODUCTION),
      .PHY_CONFIG_ENUM (PHY_CONFIG_ENUM),
      .PHY_PING_PONG_EN (PHY_PING_PONG_EN),
      .PHY_CORE_CLKS_SHARING_ENUM (PHY_CORE_CLKS_SHARING_ENUM),
      .PHY_CALIBRATED_OCT (PHY_CALIBRATED_OCT),
      .PHY_AC_CALIBRATED_OCT (PHY_AC_CALIBRATED_OCT),
      .PHY_CK_CALIBRATED_OCT (PHY_CK_CALIBRATED_OCT),
      .PHY_DATA_CALIBRATED_OCT (PHY_DATA_CALIBRATED_OCT),
      .PHY_HPS_ENABLE_EARLY_RELEASE (PHY_HPS_ENABLE_EARLY_RELEASE),
      .PLL_NUM_OF_EXTRA_CLKS (PLL_NUM_OF_EXTRA_CLKS),
      .MEM_FORMAT_ENUM (MEM_FORMAT_ENUM),
      .MEM_BURST_LENGTH (MEM_BURST_LENGTH),
      .MEM_DATA_MASK_EN (MEM_DATA_MASK_EN),
      .MEM_TTL_DATA_WIDTH (MEM_TTL_DATA_WIDTH),
      .MEM_TTL_NUM_OF_READ_GROUPS (MEM_TTL_NUM_OF_READ_GROUPS),
      .MEM_TTL_NUM_OF_WRITE_GROUPS (MEM_TTL_NUM_OF_WRITE_GROUPS),
      .DIAG_SIM_REGTEST_MODE (DIAG_SIM_REGTEST_MODE),
      .DIAG_SYNTH_FOR_SIM (DIAG_SYNTH_FOR_SIM),
      .DIAG_VERBOSE_IOAUX (DIAG_VERBOSE_IOAUX),
      .DIAG_ECLIPSE_DEBUG (DIAG_ECLIPSE_DEBUG),
      .DIAG_EXPORT_VJI (DIAG_EXPORT_VJI),
      .DIAG_INTERFACE_ID (DIAG_INTERFACE_ID),
      .DIAG_FAST_SIM (DIAG_FAST_SIM),
      .DIAG_USE_ABSTRACT_PHY (DIAG_USE_ABSTRACT_PHY),
      .SILICON_REV (SILICON_REV),
      .IS_HPS (IS_HPS),
      .IS_VID (IS_VID),
      .USER_CLK_RATIO (USER_CLK_RATIO),
      .C2P_P2C_CLK_RATIO (C2P_P2C_CLK_RATIO),
      .PHY_HMC_CLK_RATIO (PHY_HMC_CLK_RATIO),
      .DIAG_ABSTRACT_PHY_WLAT (DIAG_ABSTRACT_PHY_WLAT),
      .DIAG_ABSTRACT_PHY_RLAT (DIAG_ABSTRACT_PHY_RLAT),
      .DIAG_CPA_OUT_1_EN (DIAG_CPA_OUT_1_EN),
      .DIAG_USE_CPA_LOCK (DIAG_USE_CPA_LOCK),
      .DQS_BUS_MODE_ENUM (DQS_BUS_MODE_ENUM),
      .AC_PIN_MAP_SCHEME (AC_PIN_MAP_SCHEME),
      .NUM_OF_HMC_PORTS (NUM_OF_HMC_PORTS),
      .HMC_AVL_PROTOCOL_ENUM (HMC_AVL_PROTOCOL_ENUM),
      .HMC_CTRL_DIMM_TYPE (HMC_CTRL_DIMM_TYPE),
      .REGISTER_AFI (REGISTER_AFI),
      .SEQ_SYNTH_CPU_CLK_DIVIDE (SEQ_SYNTH_CPU_CLK_DIVIDE),
      .SEQ_SYNTH_CAL_CLK_DIVIDE (SEQ_SYNTH_CAL_CLK_DIVIDE),
      .SEQ_SIM_CPU_CLK_DIVIDE (SEQ_SIM_CPU_CLK_DIVIDE),
      .SEQ_SIM_CAL_CLK_DIVIDE (SEQ_SIM_CAL_CLK_DIVIDE),
      .SEQ_SYNTH_OSC_FREQ_MHZ (SEQ_SYNTH_OSC_FREQ_MHZ),
      .SEQ_SIM_OSC_FREQ_MHZ (SEQ_SIM_OSC_FREQ_MHZ),
      .NUM_OF_RTL_TILES (NUM_OF_RTL_TILES),
      .PRI_RDATA_TILE_INDEX (PRI_RDATA_TILE_INDEX),
      .PRI_RDATA_LANE_INDEX (PRI_RDATA_LANE_INDEX),
      .PRI_WDATA_TILE_INDEX (PRI_WDATA_TILE_INDEX),
      .PRI_WDATA_LANE_INDEX (PRI_WDATA_LANE_INDEX),
      .PRI_AC_TILE_INDEX (PRI_AC_TILE_INDEX),
      .SEC_RDATA_TILE_INDEX (SEC_RDATA_TILE_INDEX),
      .SEC_RDATA_LANE_INDEX (SEC_RDATA_LANE_INDEX),
      .SEC_WDATA_TILE_INDEX (SEC_WDATA_TILE_INDEX),
      .SEC_WDATA_LANE_INDEX (SEC_WDATA_LANE_INDEX),
      .SEC_AC_TILE_INDEX (SEC_AC_TILE_INDEX),
      .LANES_USAGE_0 (LANES_USAGE_0),
      .LANES_USAGE_1 (LANES_USAGE_1),
      .LANES_USAGE_2 (LANES_USAGE_2),
      .LANES_USAGE_3 (LANES_USAGE_3),
      .LANES_USAGE_AUTOGEN_WCNT (LANES_USAGE_AUTOGEN_WCNT),
      .PINS_USAGE_0 (PINS_USAGE_0),
      .PINS_USAGE_1 (PINS_USAGE_1),
      .PINS_USAGE_2 (PINS_USAGE_2),
      .PINS_USAGE_3 (PINS_USAGE_3),
      .PINS_USAGE_4 (PINS_USAGE_4),
      .PINS_USAGE_5 (PINS_USAGE_5),
      .PINS_USAGE_6 (PINS_USAGE_6),
      .PINS_USAGE_7 (PINS_USAGE_7),
      .PINS_USAGE_8 (PINS_USAGE_8),
      .PINS_USAGE_9 (PINS_USAGE_9),
      .PINS_USAGE_10 (PINS_USAGE_10),
      .PINS_USAGE_11 (PINS_USAGE_11),
      .PINS_USAGE_12 (PINS_USAGE_12),
      .PINS_USAGE_AUTOGEN_WCNT (PINS_USAGE_AUTOGEN_WCNT),
      .PINS_RATE_0 (PINS_RATE_0),
      .PINS_RATE_1 (PINS_RATE_1),
      .PINS_RATE_2 (PINS_RATE_2),
      .PINS_RATE_3 (PINS_RATE_3),
      .PINS_RATE_4 (PINS_RATE_4),
      .PINS_RATE_5 (PINS_RATE_5),
      .PINS_RATE_6 (PINS_RATE_6),
      .PINS_RATE_7 (PINS_RATE_7),
      .PINS_RATE_8 (PINS_RATE_8),
      .PINS_RATE_9 (PINS_RATE_9),
      .PINS_RATE_10 (PINS_RATE_10),
      .PINS_RATE_11 (PINS_RATE_11),
      .PINS_RATE_12 (PINS_RATE_12),
      .PINS_RATE_AUTOGEN_WCNT (PINS_RATE_AUTOGEN_WCNT),
      .PINS_WDB_0 (PINS_WDB_0),
      .PINS_WDB_1 (PINS_WDB_1),
      .PINS_WDB_2 (PINS_WDB_2),
      .PINS_WDB_3 (PINS_WDB_3),
      .PINS_WDB_4 (PINS_WDB_4),
      .PINS_WDB_5 (PINS_WDB_5),
      .PINS_WDB_6 (PINS_WDB_6),
      .PINS_WDB_7 (PINS_WDB_7),
      .PINS_WDB_8 (PINS_WDB_8),
      .PINS_WDB_9 (PINS_WDB_9),
      .PINS_WDB_10 (PINS_WDB_10),
      .PINS_WDB_11 (PINS_WDB_11),
      .PINS_WDB_12 (PINS_WDB_12),
      .PINS_WDB_13 (PINS_WDB_13),
      .PINS_WDB_14 (PINS_WDB_14),
      .PINS_WDB_15 (PINS_WDB_15),
      .PINS_WDB_16 (PINS_WDB_16),
      .PINS_WDB_17 (PINS_WDB_17),
      .PINS_WDB_18 (PINS_WDB_18),
      .PINS_WDB_19 (PINS_WDB_19),
      .PINS_WDB_20 (PINS_WDB_20),
      .PINS_WDB_21 (PINS_WDB_21),
      .PINS_WDB_22 (PINS_WDB_22),
      .PINS_WDB_23 (PINS_WDB_23),
      .PINS_WDB_24 (PINS_WDB_24),
      .PINS_WDB_25 (PINS_WDB_25),
      .PINS_WDB_26 (PINS_WDB_26),
      .PINS_WDB_27 (PINS_WDB_27),
      .PINS_WDB_28 (PINS_WDB_28),
      .PINS_WDB_29 (PINS_WDB_29),
      .PINS_WDB_30 (PINS_WDB_30),
      .PINS_WDB_31 (PINS_WDB_31),
      .PINS_WDB_32 (PINS_WDB_32),
      .PINS_WDB_33 (PINS_WDB_33),
      .PINS_WDB_34 (PINS_WDB_34),
      .PINS_WDB_35 (PINS_WDB_35),
      .PINS_WDB_36 (PINS_WDB_36),
      .PINS_WDB_37 (PINS_WDB_37),
      .PINS_WDB_38 (PINS_WDB_38),
      .PINS_WDB_AUTOGEN_WCNT (PINS_WDB_AUTOGEN_WCNT),
      .PINS_DATA_IN_MODE_0 (PINS_DATA_IN_MODE_0),
      .PINS_DATA_IN_MODE_1 (PINS_DATA_IN_MODE_1),
      .PINS_DATA_IN_MODE_2 (PINS_DATA_IN_MODE_2),
      .PINS_DATA_IN_MODE_3 (PINS_DATA_IN_MODE_3),
      .PINS_DATA_IN_MODE_4 (PINS_DATA_IN_MODE_4),
      .PINS_DATA_IN_MODE_5 (PINS_DATA_IN_MODE_5),
      .PINS_DATA_IN_MODE_6 (PINS_DATA_IN_MODE_6),
      .PINS_DATA_IN_MODE_7 (PINS_DATA_IN_MODE_7),
      .PINS_DATA_IN_MODE_8 (PINS_DATA_IN_MODE_8),
      .PINS_DATA_IN_MODE_9 (PINS_DATA_IN_MODE_9),
      .PINS_DATA_IN_MODE_10 (PINS_DATA_IN_MODE_10),
      .PINS_DATA_IN_MODE_11 (PINS_DATA_IN_MODE_11),
      .PINS_DATA_IN_MODE_12 (PINS_DATA_IN_MODE_12),
      .PINS_DATA_IN_MODE_13 (PINS_DATA_IN_MODE_13),
      .PINS_DATA_IN_MODE_14 (PINS_DATA_IN_MODE_14),
      .PINS_DATA_IN_MODE_15 (PINS_DATA_IN_MODE_15),
      .PINS_DATA_IN_MODE_16 (PINS_DATA_IN_MODE_16),
      .PINS_DATA_IN_MODE_17 (PINS_DATA_IN_MODE_17),
      .PINS_DATA_IN_MODE_18 (PINS_DATA_IN_MODE_18),
      .PINS_DATA_IN_MODE_19 (PINS_DATA_IN_MODE_19),
      .PINS_DATA_IN_MODE_20 (PINS_DATA_IN_MODE_20),
      .PINS_DATA_IN_MODE_21 (PINS_DATA_IN_MODE_21),
      .PINS_DATA_IN_MODE_22 (PINS_DATA_IN_MODE_22),
      .PINS_DATA_IN_MODE_23 (PINS_DATA_IN_MODE_23),
      .PINS_DATA_IN_MODE_24 (PINS_DATA_IN_MODE_24),
      .PINS_DATA_IN_MODE_25 (PINS_DATA_IN_MODE_25),
      .PINS_DATA_IN_MODE_26 (PINS_DATA_IN_MODE_26),
      .PINS_DATA_IN_MODE_27 (PINS_DATA_IN_MODE_27),
      .PINS_DATA_IN_MODE_28 (PINS_DATA_IN_MODE_28),
      .PINS_DATA_IN_MODE_29 (PINS_DATA_IN_MODE_29),
      .PINS_DATA_IN_MODE_30 (PINS_DATA_IN_MODE_30),
      .PINS_DATA_IN_MODE_31 (PINS_DATA_IN_MODE_31),
      .PINS_DATA_IN_MODE_32 (PINS_DATA_IN_MODE_32),
      .PINS_DATA_IN_MODE_33 (PINS_DATA_IN_MODE_33),
      .PINS_DATA_IN_MODE_34 (PINS_DATA_IN_MODE_34),
      .PINS_DATA_IN_MODE_35 (PINS_DATA_IN_MODE_35),
      .PINS_DATA_IN_MODE_36 (PINS_DATA_IN_MODE_36),
      .PINS_DATA_IN_MODE_37 (PINS_DATA_IN_MODE_37),
      .PINS_DATA_IN_MODE_38 (PINS_DATA_IN_MODE_38),
      .PINS_DATA_IN_MODE_AUTOGEN_WCNT (PINS_DATA_IN_MODE_AUTOGEN_WCNT),
      .PINS_C2L_DRIVEN_0 (PINS_C2L_DRIVEN_0),
      .PINS_C2L_DRIVEN_1 (PINS_C2L_DRIVEN_1),
      .PINS_C2L_DRIVEN_2 (PINS_C2L_DRIVEN_2),
      .PINS_C2L_DRIVEN_3 (PINS_C2L_DRIVEN_3),
      .PINS_C2L_DRIVEN_4 (PINS_C2L_DRIVEN_4),
      .PINS_C2L_DRIVEN_5 (PINS_C2L_DRIVEN_5),
      .PINS_C2L_DRIVEN_6 (PINS_C2L_DRIVEN_6),
      .PINS_C2L_DRIVEN_7 (PINS_C2L_DRIVEN_7),
      .PINS_C2L_DRIVEN_8 (PINS_C2L_DRIVEN_8),
      .PINS_C2L_DRIVEN_9 (PINS_C2L_DRIVEN_9),
      .PINS_C2L_DRIVEN_10 (PINS_C2L_DRIVEN_10),
      .PINS_C2L_DRIVEN_11 (PINS_C2L_DRIVEN_11),
      .PINS_C2L_DRIVEN_12 (PINS_C2L_DRIVEN_12),
      .PINS_C2L_DRIVEN_AUTOGEN_WCNT (PINS_C2L_DRIVEN_AUTOGEN_WCNT),
      .PINS_DB_IN_BYPASS_0 (PINS_DB_IN_BYPASS_0),
      .PINS_DB_IN_BYPASS_1 (PINS_DB_IN_BYPASS_1),
      .PINS_DB_IN_BYPASS_2 (PINS_DB_IN_BYPASS_2),
      .PINS_DB_IN_BYPASS_3 (PINS_DB_IN_BYPASS_3),
      .PINS_DB_IN_BYPASS_4 (PINS_DB_IN_BYPASS_4),
      .PINS_DB_IN_BYPASS_5 (PINS_DB_IN_BYPASS_5),
      .PINS_DB_IN_BYPASS_6 (PINS_DB_IN_BYPASS_6),
      .PINS_DB_IN_BYPASS_7 (PINS_DB_IN_BYPASS_7),
      .PINS_DB_IN_BYPASS_8 (PINS_DB_IN_BYPASS_8),
      .PINS_DB_IN_BYPASS_9 (PINS_DB_IN_BYPASS_9),
      .PINS_DB_IN_BYPASS_10 (PINS_DB_IN_BYPASS_10),
      .PINS_DB_IN_BYPASS_11 (PINS_DB_IN_BYPASS_11),
      .PINS_DB_IN_BYPASS_12 (PINS_DB_IN_BYPASS_12),
      .PINS_DB_IN_BYPASS_AUTOGEN_WCNT (PINS_DB_IN_BYPASS_AUTOGEN_WCNT),
      .PINS_DB_OUT_BYPASS_0 (PINS_DB_OUT_BYPASS_0),
      .PINS_DB_OUT_BYPASS_1 (PINS_DB_OUT_BYPASS_1),
      .PINS_DB_OUT_BYPASS_2 (PINS_DB_OUT_BYPASS_2),
      .PINS_DB_OUT_BYPASS_3 (PINS_DB_OUT_BYPASS_3),
      .PINS_DB_OUT_BYPASS_4 (PINS_DB_OUT_BYPASS_4),
      .PINS_DB_OUT_BYPASS_5 (PINS_DB_OUT_BYPASS_5),
      .PINS_DB_OUT_BYPASS_6 (PINS_DB_OUT_BYPASS_6),
      .PINS_DB_OUT_BYPASS_7 (PINS_DB_OUT_BYPASS_7),
      .PINS_DB_OUT_BYPASS_8 (PINS_DB_OUT_BYPASS_8),
      .PINS_DB_OUT_BYPASS_9 (PINS_DB_OUT_BYPASS_9),
      .PINS_DB_OUT_BYPASS_10 (PINS_DB_OUT_BYPASS_10),
      .PINS_DB_OUT_BYPASS_11 (PINS_DB_OUT_BYPASS_11),
      .PINS_DB_OUT_BYPASS_12 (PINS_DB_OUT_BYPASS_12),
      .PINS_DB_OUT_BYPASS_AUTOGEN_WCNT (PINS_DB_OUT_BYPASS_AUTOGEN_WCNT),
      .PINS_DB_OE_BYPASS_0 (PINS_DB_OE_BYPASS_0),
      .PINS_DB_OE_BYPASS_1 (PINS_DB_OE_BYPASS_1),
      .PINS_DB_OE_BYPASS_2 (PINS_DB_OE_BYPASS_2),
      .PINS_DB_OE_BYPASS_3 (PINS_DB_OE_BYPASS_3),
      .PINS_DB_OE_BYPASS_4 (PINS_DB_OE_BYPASS_4),
      .PINS_DB_OE_BYPASS_5 (PINS_DB_OE_BYPASS_5),
      .PINS_DB_OE_BYPASS_6 (PINS_DB_OE_BYPASS_6),
      .PINS_DB_OE_BYPASS_7 (PINS_DB_OE_BYPASS_7),
      .PINS_DB_OE_BYPASS_8 (PINS_DB_OE_BYPASS_8),
      .PINS_DB_OE_BYPASS_9 (PINS_DB_OE_BYPASS_9),
      .PINS_DB_OE_BYPASS_10 (PINS_DB_OE_BYPASS_10),
      .PINS_DB_OE_BYPASS_11 (PINS_DB_OE_BYPASS_11),
      .PINS_DB_OE_BYPASS_12 (PINS_DB_OE_BYPASS_12),
      .PINS_DB_OE_BYPASS_AUTOGEN_WCNT (PINS_DB_OE_BYPASS_AUTOGEN_WCNT),
      .PINS_INVERT_WR_0 (PINS_INVERT_WR_0),
      .PINS_INVERT_WR_1 (PINS_INVERT_WR_1),
      .PINS_INVERT_WR_2 (PINS_INVERT_WR_2),
      .PINS_INVERT_WR_3 (PINS_INVERT_WR_3),
      .PINS_INVERT_WR_4 (PINS_INVERT_WR_4),
      .PINS_INVERT_WR_5 (PINS_INVERT_WR_5),
      .PINS_INVERT_WR_6 (PINS_INVERT_WR_6),
      .PINS_INVERT_WR_7 (PINS_INVERT_WR_7),
      .PINS_INVERT_WR_8 (PINS_INVERT_WR_8),
      .PINS_INVERT_WR_9 (PINS_INVERT_WR_9),
      .PINS_INVERT_WR_10 (PINS_INVERT_WR_10),
      .PINS_INVERT_WR_11 (PINS_INVERT_WR_11),
      .PINS_INVERT_WR_12 (PINS_INVERT_WR_12),
      .PINS_INVERT_WR_AUTOGEN_WCNT (PINS_INVERT_WR_AUTOGEN_WCNT),
      .PINS_INVERT_OE_0 (PINS_INVERT_OE_0),
      .PINS_INVERT_OE_1 (PINS_INVERT_OE_1),
      .PINS_INVERT_OE_2 (PINS_INVERT_OE_2),
      .PINS_INVERT_OE_3 (PINS_INVERT_OE_3),
      .PINS_INVERT_OE_4 (PINS_INVERT_OE_4),
      .PINS_INVERT_OE_5 (PINS_INVERT_OE_5),
      .PINS_INVERT_OE_6 (PINS_INVERT_OE_6),
      .PINS_INVERT_OE_7 (PINS_INVERT_OE_7),
      .PINS_INVERT_OE_8 (PINS_INVERT_OE_8),
      .PINS_INVERT_OE_9 (PINS_INVERT_OE_9),
      .PINS_INVERT_OE_10 (PINS_INVERT_OE_10),
      .PINS_INVERT_OE_11 (PINS_INVERT_OE_11),
      .PINS_INVERT_OE_12 (PINS_INVERT_OE_12),
      .PINS_INVERT_OE_AUTOGEN_WCNT (PINS_INVERT_OE_AUTOGEN_WCNT),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_0 (PINS_AC_HMC_DATA_OVERRIDE_ENA_0),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_1 (PINS_AC_HMC_DATA_OVERRIDE_ENA_1),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_2 (PINS_AC_HMC_DATA_OVERRIDE_ENA_2),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_3 (PINS_AC_HMC_DATA_OVERRIDE_ENA_3),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_4 (PINS_AC_HMC_DATA_OVERRIDE_ENA_4),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_5 (PINS_AC_HMC_DATA_OVERRIDE_ENA_5),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_6 (PINS_AC_HMC_DATA_OVERRIDE_ENA_6),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_7 (PINS_AC_HMC_DATA_OVERRIDE_ENA_7),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_8 (PINS_AC_HMC_DATA_OVERRIDE_ENA_8),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_9 (PINS_AC_HMC_DATA_OVERRIDE_ENA_9),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_10 (PINS_AC_HMC_DATA_OVERRIDE_ENA_10),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_11 (PINS_AC_HMC_DATA_OVERRIDE_ENA_11),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_12 (PINS_AC_HMC_DATA_OVERRIDE_ENA_12),
      .PINS_AC_HMC_DATA_OVERRIDE_ENA_AUTOGEN_WCNT (PINS_AC_HMC_DATA_OVERRIDE_ENA_AUTOGEN_WCNT),
      .PINS_OCT_MODE_0 (PINS_OCT_MODE_0),
      .PINS_OCT_MODE_1 (PINS_OCT_MODE_1),
      .PINS_OCT_MODE_2 (PINS_OCT_MODE_2),
      .PINS_OCT_MODE_3 (PINS_OCT_MODE_3),
      .PINS_OCT_MODE_4 (PINS_OCT_MODE_4),
      .PINS_OCT_MODE_5 (PINS_OCT_MODE_5),
      .PINS_OCT_MODE_6 (PINS_OCT_MODE_6),
      .PINS_OCT_MODE_7 (PINS_OCT_MODE_7),
      .PINS_OCT_MODE_8 (PINS_OCT_MODE_8),
      .PINS_OCT_MODE_9 (PINS_OCT_MODE_9),
      .PINS_OCT_MODE_10 (PINS_OCT_MODE_10),
      .PINS_OCT_MODE_11 (PINS_OCT_MODE_11),
      .PINS_OCT_MODE_12 (PINS_OCT_MODE_12),
      .PINS_OCT_MODE_AUTOGEN_WCNT (PINS_OCT_MODE_AUTOGEN_WCNT),
      .PINS_GPIO_MODE_0 (PINS_GPIO_MODE_0),
      .PINS_GPIO_MODE_1 (PINS_GPIO_MODE_1),
      .PINS_GPIO_MODE_2 (PINS_GPIO_MODE_2),
      .PINS_GPIO_MODE_3 (PINS_GPIO_MODE_3),
      .PINS_GPIO_MODE_4 (PINS_GPIO_MODE_4),
      .PINS_GPIO_MODE_5 (PINS_GPIO_MODE_5),
      .PINS_GPIO_MODE_6 (PINS_GPIO_MODE_6),
      .PINS_GPIO_MODE_7 (PINS_GPIO_MODE_7),
      .PINS_GPIO_MODE_8 (PINS_GPIO_MODE_8),
      .PINS_GPIO_MODE_9 (PINS_GPIO_MODE_9),
      .PINS_GPIO_MODE_10 (PINS_GPIO_MODE_10),
      .PINS_GPIO_MODE_11 (PINS_GPIO_MODE_11),
      .PINS_GPIO_MODE_12 (PINS_GPIO_MODE_12),
      .PINS_GPIO_MODE_AUTOGEN_WCNT (PINS_GPIO_MODE_AUTOGEN_WCNT),
      .UNUSED_MEM_PINS_PINLOC_0 (UNUSED_MEM_PINS_PINLOC_0),
      .UNUSED_MEM_PINS_PINLOC_1 (UNUSED_MEM_PINS_PINLOC_1),
      .UNUSED_MEM_PINS_PINLOC_2 (UNUSED_MEM_PINS_PINLOC_2),
      .UNUSED_MEM_PINS_PINLOC_3 (UNUSED_MEM_PINS_PINLOC_3),
      .UNUSED_MEM_PINS_PINLOC_4 (UNUSED_MEM_PINS_PINLOC_4),
      .UNUSED_MEM_PINS_PINLOC_5 (UNUSED_MEM_PINS_PINLOC_5),
      .UNUSED_MEM_PINS_PINLOC_6 (UNUSED_MEM_PINS_PINLOC_6),
      .UNUSED_MEM_PINS_PINLOC_7 (UNUSED_MEM_PINS_PINLOC_7),
      .UNUSED_MEM_PINS_PINLOC_8 (UNUSED_MEM_PINS_PINLOC_8),
      .UNUSED_MEM_PINS_PINLOC_9 (UNUSED_MEM_PINS_PINLOC_9),
      .UNUSED_MEM_PINS_PINLOC_10 (UNUSED_MEM_PINS_PINLOC_10),
      .UNUSED_MEM_PINS_PINLOC_11 (UNUSED_MEM_PINS_PINLOC_11),
      .UNUSED_MEM_PINS_PINLOC_12 (UNUSED_MEM_PINS_PINLOC_12),
      .UNUSED_MEM_PINS_PINLOC_13 (UNUSED_MEM_PINS_PINLOC_13),
      .UNUSED_MEM_PINS_PINLOC_14 (UNUSED_MEM_PINS_PINLOC_14),
      .UNUSED_MEM_PINS_PINLOC_15 (UNUSED_MEM_PINS_PINLOC_15),
      .UNUSED_MEM_PINS_PINLOC_16 (UNUSED_MEM_PINS_PINLOC_16),
      .UNUSED_MEM_PINS_PINLOC_17 (UNUSED_MEM_PINS_PINLOC_17),
      .UNUSED_MEM_PINS_PINLOC_18 (UNUSED_MEM_PINS_PINLOC_18),
      .UNUSED_MEM_PINS_PINLOC_19 (UNUSED_MEM_PINS_PINLOC_19),
      .UNUSED_MEM_PINS_PINLOC_20 (UNUSED_MEM_PINS_PINLOC_20),
      .UNUSED_MEM_PINS_PINLOC_21 (UNUSED_MEM_PINS_PINLOC_21),
      .UNUSED_MEM_PINS_PINLOC_22 (UNUSED_MEM_PINS_PINLOC_22),
      .UNUSED_MEM_PINS_PINLOC_23 (UNUSED_MEM_PINS_PINLOC_23),
      .UNUSED_MEM_PINS_PINLOC_24 (UNUSED_MEM_PINS_PINLOC_24),
      .UNUSED_MEM_PINS_PINLOC_25 (UNUSED_MEM_PINS_PINLOC_25),
      .UNUSED_MEM_PINS_PINLOC_26 (UNUSED_MEM_PINS_PINLOC_26),
      .UNUSED_MEM_PINS_PINLOC_27 (UNUSED_MEM_PINS_PINLOC_27),
      .UNUSED_MEM_PINS_PINLOC_28 (UNUSED_MEM_PINS_PINLOC_28),
      .UNUSED_MEM_PINS_PINLOC_29 (UNUSED_MEM_PINS_PINLOC_29),
      .UNUSED_MEM_PINS_PINLOC_30 (UNUSED_MEM_PINS_PINLOC_30),
      .UNUSED_MEM_PINS_PINLOC_31 (UNUSED_MEM_PINS_PINLOC_31),
      .UNUSED_MEM_PINS_PINLOC_32 (UNUSED_MEM_PINS_PINLOC_32),
      .UNUSED_MEM_PINS_PINLOC_33 (UNUSED_MEM_PINS_PINLOC_33),
      .UNUSED_MEM_PINS_PINLOC_34 (UNUSED_MEM_PINS_PINLOC_34),
      .UNUSED_MEM_PINS_PINLOC_35 (UNUSED_MEM_PINS_PINLOC_35),
      .UNUSED_MEM_PINS_PINLOC_36 (UNUSED_MEM_PINS_PINLOC_36),
      .UNUSED_MEM_PINS_PINLOC_37 (UNUSED_MEM_PINS_PINLOC_37),
      .UNUSED_MEM_PINS_PINLOC_38 (UNUSED_MEM_PINS_PINLOC_38),
      .UNUSED_MEM_PINS_PINLOC_39 (UNUSED_MEM_PINS_PINLOC_39),
      .UNUSED_MEM_PINS_PINLOC_40 (UNUSED_MEM_PINS_PINLOC_40),
      .UNUSED_MEM_PINS_PINLOC_41 (UNUSED_MEM_PINS_PINLOC_41),
      .UNUSED_MEM_PINS_PINLOC_42 (UNUSED_MEM_PINS_PINLOC_42),
      .UNUSED_MEM_PINS_PINLOC_43 (UNUSED_MEM_PINS_PINLOC_43),
      .UNUSED_MEM_PINS_PINLOC_44 (UNUSED_MEM_PINS_PINLOC_44),
      .UNUSED_MEM_PINS_PINLOC_45 (UNUSED_MEM_PINS_PINLOC_45),
      .UNUSED_MEM_PINS_PINLOC_46 (UNUSED_MEM_PINS_PINLOC_46),
      .UNUSED_MEM_PINS_PINLOC_47 (UNUSED_MEM_PINS_PINLOC_47),
      .UNUSED_MEM_PINS_PINLOC_48 (UNUSED_MEM_PINS_PINLOC_48),
      .UNUSED_MEM_PINS_PINLOC_49 (UNUSED_MEM_PINS_PINLOC_49),
      .UNUSED_MEM_PINS_PINLOC_50 (UNUSED_MEM_PINS_PINLOC_50),
      .UNUSED_MEM_PINS_PINLOC_51 (UNUSED_MEM_PINS_PINLOC_51),
      .UNUSED_MEM_PINS_PINLOC_52 (UNUSED_MEM_PINS_PINLOC_52),
      .UNUSED_MEM_PINS_PINLOC_53 (UNUSED_MEM_PINS_PINLOC_53),
      .UNUSED_MEM_PINS_PINLOC_54 (UNUSED_MEM_PINS_PINLOC_54),
      .UNUSED_MEM_PINS_PINLOC_55 (UNUSED_MEM_PINS_PINLOC_55),
      .UNUSED_MEM_PINS_PINLOC_56 (UNUSED_MEM_PINS_PINLOC_56),
      .UNUSED_MEM_PINS_PINLOC_57 (UNUSED_MEM_PINS_PINLOC_57),
      .UNUSED_MEM_PINS_PINLOC_58 (UNUSED_MEM_PINS_PINLOC_58),
      .UNUSED_MEM_PINS_PINLOC_59 (UNUSED_MEM_PINS_PINLOC_59),
      .UNUSED_MEM_PINS_PINLOC_60 (UNUSED_MEM_PINS_PINLOC_60),
      .UNUSED_MEM_PINS_PINLOC_61 (UNUSED_MEM_PINS_PINLOC_61),
      .UNUSED_MEM_PINS_PINLOC_62 (UNUSED_MEM_PINS_PINLOC_62),
      .UNUSED_MEM_PINS_PINLOC_63 (UNUSED_MEM_PINS_PINLOC_63),
      .UNUSED_MEM_PINS_PINLOC_64 (UNUSED_MEM_PINS_PINLOC_64),
      .UNUSED_MEM_PINS_PINLOC_65 (UNUSED_MEM_PINS_PINLOC_65),
      .UNUSED_MEM_PINS_PINLOC_66 (UNUSED_MEM_PINS_PINLOC_66),
      .UNUSED_MEM_PINS_PINLOC_67 (UNUSED_MEM_PINS_PINLOC_67),
      .UNUSED_MEM_PINS_PINLOC_68 (UNUSED_MEM_PINS_PINLOC_68),
      .UNUSED_MEM_PINS_PINLOC_69 (UNUSED_MEM_PINS_PINLOC_69),
      .UNUSED_MEM_PINS_PINLOC_70 (UNUSED_MEM_PINS_PINLOC_70),
      .UNUSED_MEM_PINS_PINLOC_71 (UNUSED_MEM_PINS_PINLOC_71),
      .UNUSED_MEM_PINS_PINLOC_72 (UNUSED_MEM_PINS_PINLOC_72),
      .UNUSED_MEM_PINS_PINLOC_73 (UNUSED_MEM_PINS_PINLOC_73),
      .UNUSED_MEM_PINS_PINLOC_74 (UNUSED_MEM_PINS_PINLOC_74),
      .UNUSED_MEM_PINS_PINLOC_75 (UNUSED_MEM_PINS_PINLOC_75),
      .UNUSED_MEM_PINS_PINLOC_76 (UNUSED_MEM_PINS_PINLOC_76),
      .UNUSED_MEM_PINS_PINLOC_77 (UNUSED_MEM_PINS_PINLOC_77),
      .UNUSED_MEM_PINS_PINLOC_78 (UNUSED_MEM_PINS_PINLOC_78),
      .UNUSED_MEM_PINS_PINLOC_79 (UNUSED_MEM_PINS_PINLOC_79),
      .UNUSED_MEM_PINS_PINLOC_80 (UNUSED_MEM_PINS_PINLOC_80),
      .UNUSED_MEM_PINS_PINLOC_81 (UNUSED_MEM_PINS_PINLOC_81),
      .UNUSED_MEM_PINS_PINLOC_82 (UNUSED_MEM_PINS_PINLOC_82),
      .UNUSED_MEM_PINS_PINLOC_83 (UNUSED_MEM_PINS_PINLOC_83),
      .UNUSED_MEM_PINS_PINLOC_84 (UNUSED_MEM_PINS_PINLOC_84),
      .UNUSED_MEM_PINS_PINLOC_85 (UNUSED_MEM_PINS_PINLOC_85),
      .UNUSED_MEM_PINS_PINLOC_86 (UNUSED_MEM_PINS_PINLOC_86),
      .UNUSED_MEM_PINS_PINLOC_87 (UNUSED_MEM_PINS_PINLOC_87),
      .UNUSED_MEM_PINS_PINLOC_88 (UNUSED_MEM_PINS_PINLOC_88),
      .UNUSED_MEM_PINS_PINLOC_89 (UNUSED_MEM_PINS_PINLOC_89),
      .UNUSED_MEM_PINS_PINLOC_90 (UNUSED_MEM_PINS_PINLOC_90),
      .UNUSED_MEM_PINS_PINLOC_91 (UNUSED_MEM_PINS_PINLOC_91),
      .UNUSED_MEM_PINS_PINLOC_92 (UNUSED_MEM_PINS_PINLOC_92),
      .UNUSED_MEM_PINS_PINLOC_93 (UNUSED_MEM_PINS_PINLOC_93),
      .UNUSED_MEM_PINS_PINLOC_94 (UNUSED_MEM_PINS_PINLOC_94),
      .UNUSED_MEM_PINS_PINLOC_95 (UNUSED_MEM_PINS_PINLOC_95),
      .UNUSED_MEM_PINS_PINLOC_96 (UNUSED_MEM_PINS_PINLOC_96),
      .UNUSED_MEM_PINS_PINLOC_97 (UNUSED_MEM_PINS_PINLOC_97),
      .UNUSED_MEM_PINS_PINLOC_98 (UNUSED_MEM_PINS_PINLOC_98),
      .UNUSED_MEM_PINS_PINLOC_99 (UNUSED_MEM_PINS_PINLOC_99),
      .UNUSED_MEM_PINS_PINLOC_100 (UNUSED_MEM_PINS_PINLOC_100),
      .UNUSED_MEM_PINS_PINLOC_101 (UNUSED_MEM_PINS_PINLOC_101),
      .UNUSED_MEM_PINS_PINLOC_102 (UNUSED_MEM_PINS_PINLOC_102),
      .UNUSED_MEM_PINS_PINLOC_103 (UNUSED_MEM_PINS_PINLOC_103),
      .UNUSED_MEM_PINS_PINLOC_104 (UNUSED_MEM_PINS_PINLOC_104),
      .UNUSED_MEM_PINS_PINLOC_105 (UNUSED_MEM_PINS_PINLOC_105),
      .UNUSED_MEM_PINS_PINLOC_106 (UNUSED_MEM_PINS_PINLOC_106),
      .UNUSED_MEM_PINS_PINLOC_107 (UNUSED_MEM_PINS_PINLOC_107),
      .UNUSED_MEM_PINS_PINLOC_108 (UNUSED_MEM_PINS_PINLOC_108),
      .UNUSED_MEM_PINS_PINLOC_109 (UNUSED_MEM_PINS_PINLOC_109),
      .UNUSED_MEM_PINS_PINLOC_110 (UNUSED_MEM_PINS_PINLOC_110),
      .UNUSED_MEM_PINS_PINLOC_111 (UNUSED_MEM_PINS_PINLOC_111),
      .UNUSED_MEM_PINS_PINLOC_112 (UNUSED_MEM_PINS_PINLOC_112),
      .UNUSED_MEM_PINS_PINLOC_113 (UNUSED_MEM_PINS_PINLOC_113),
      .UNUSED_MEM_PINS_PINLOC_114 (UNUSED_MEM_PINS_PINLOC_114),
      .UNUSED_MEM_PINS_PINLOC_115 (UNUSED_MEM_PINS_PINLOC_115),
      .UNUSED_MEM_PINS_PINLOC_116 (UNUSED_MEM_PINS_PINLOC_116),
      .UNUSED_MEM_PINS_PINLOC_117 (UNUSED_MEM_PINS_PINLOC_117),
      .UNUSED_MEM_PINS_PINLOC_118 (UNUSED_MEM_PINS_PINLOC_118),
      .UNUSED_MEM_PINS_PINLOC_119 (UNUSED_MEM_PINS_PINLOC_119),
      .UNUSED_MEM_PINS_PINLOC_120 (UNUSED_MEM_PINS_PINLOC_120),
      .UNUSED_MEM_PINS_PINLOC_121 (UNUSED_MEM_PINS_PINLOC_121),
      .UNUSED_MEM_PINS_PINLOC_122 (UNUSED_MEM_PINS_PINLOC_122),
      .UNUSED_MEM_PINS_PINLOC_123 (UNUSED_MEM_PINS_PINLOC_123),
      .UNUSED_MEM_PINS_PINLOC_124 (UNUSED_MEM_PINS_PINLOC_124),
      .UNUSED_MEM_PINS_PINLOC_125 (UNUSED_MEM_PINS_PINLOC_125),
      .UNUSED_MEM_PINS_PINLOC_126 (UNUSED_MEM_PINS_PINLOC_126),
      .UNUSED_MEM_PINS_PINLOC_127 (UNUSED_MEM_PINS_PINLOC_127),
      .UNUSED_MEM_PINS_PINLOC_128 (UNUSED_MEM_PINS_PINLOC_128),
      .UNUSED_MEM_PINS_PINLOC_AUTOGEN_WCNT (UNUSED_MEM_PINS_PINLOC_AUTOGEN_WCNT),
      .UNUSED_DQS_BUSES_LANELOC_0 (UNUSED_DQS_BUSES_LANELOC_0),
      .UNUSED_DQS_BUSES_LANELOC_1 (UNUSED_DQS_BUSES_LANELOC_1),
      .UNUSED_DQS_BUSES_LANELOC_2 (UNUSED_DQS_BUSES_LANELOC_2),
      .UNUSED_DQS_BUSES_LANELOC_3 (UNUSED_DQS_BUSES_LANELOC_3),
      .UNUSED_DQS_BUSES_LANELOC_4 (UNUSED_DQS_BUSES_LANELOC_4),
      .UNUSED_DQS_BUSES_LANELOC_5 (UNUSED_DQS_BUSES_LANELOC_5),
      .UNUSED_DQS_BUSES_LANELOC_6 (UNUSED_DQS_BUSES_LANELOC_6),
      .UNUSED_DQS_BUSES_LANELOC_7 (UNUSED_DQS_BUSES_LANELOC_7),
      .UNUSED_DQS_BUSES_LANELOC_8 (UNUSED_DQS_BUSES_LANELOC_8),
      .UNUSED_DQS_BUSES_LANELOC_9 (UNUSED_DQS_BUSES_LANELOC_9),
      .UNUSED_DQS_BUSES_LANELOC_10 (UNUSED_DQS_BUSES_LANELOC_10),
      .UNUSED_DQS_BUSES_LANELOC_AUTOGEN_WCNT (UNUSED_DQS_BUSES_LANELOC_AUTOGEN_WCNT),
      .CENTER_TIDS_0 (CENTER_TIDS_0),
      .CENTER_TIDS_1 (CENTER_TIDS_1),
      .CENTER_TIDS_2 (CENTER_TIDS_2),
      .CENTER_TIDS_AUTOGEN_WCNT (CENTER_TIDS_AUTOGEN_WCNT),
      .HMC_TIDS_0 (HMC_TIDS_0),
      .HMC_TIDS_1 (HMC_TIDS_1),
      .HMC_TIDS_2 (HMC_TIDS_2),
      .HMC_TIDS_AUTOGEN_WCNT (HMC_TIDS_AUTOGEN_WCNT),
      .LANE_TIDS_0 (LANE_TIDS_0),
      .LANE_TIDS_1 (LANE_TIDS_1),
      .LANE_TIDS_2 (LANE_TIDS_2),
      .LANE_TIDS_3 (LANE_TIDS_3),
      .LANE_TIDS_4 (LANE_TIDS_4),
      .LANE_TIDS_5 (LANE_TIDS_5),
      .LANE_TIDS_6 (LANE_TIDS_6),
      .LANE_TIDS_7 (LANE_TIDS_7),
      .LANE_TIDS_8 (LANE_TIDS_8),
      .LANE_TIDS_9 (LANE_TIDS_9),
      .LANE_TIDS_AUTOGEN_WCNT (LANE_TIDS_AUTOGEN_WCNT),
      .PREAMBLE_MODE (PREAMBLE_MODE),
      .DBI_WR_ENABLE (DBI_WR_ENABLE),
      .DBI_RD_ENABLE (DBI_RD_ENABLE),
      .CRC_EN (CRC_EN),
      .SWAP_DQS_A_B (SWAP_DQS_A_B),
      .DQS_PACK_MODE (DQS_PACK_MODE),
      .OCT_SIZE (OCT_SIZE),
      .DBC_WB_RESERVED_ENTRY (DBC_WB_RESERVED_ENTRY),
      .DLL_MODE (DLL_MODE),
      .DLL_CODEWORD (DLL_CODEWORD),
      .ABPHY_WRITE_PROTOCOL (ABPHY_WRITE_PROTOCOL),
      .PHY_USERMODE_OCT (PHY_USERMODE_OCT),
      .PHY_PERIODIC_OCT_RECAL (PHY_PERIODIC_OCT_RECAL),
      .PHY_HAS_DCC (PHY_HAS_DCC),
      .PRI_HMC_CFG_ENABLE_ECC (PRI_HMC_CFG_ENABLE_ECC),
      .PRI_HMC_CFG_REORDER_DATA (PRI_HMC_CFG_REORDER_DATA),
      .PRI_HMC_CFG_REORDER_READ (PRI_HMC_CFG_REORDER_READ),
      .PRI_HMC_CFG_REORDER_RDATA (PRI_HMC_CFG_REORDER_RDATA),
      .PRI_HMC_CFG_STARVE_LIMIT (PRI_HMC_CFG_STARVE_LIMIT),
      .PRI_HMC_CFG_DQS_TRACKING_EN (PRI_HMC_CFG_DQS_TRACKING_EN),
      .PRI_HMC_CFG_ARBITER_TYPE (PRI_HMC_CFG_ARBITER_TYPE),
      .PRI_HMC_CFG_OPEN_PAGE_EN (PRI_HMC_CFG_OPEN_PAGE_EN),
      .PRI_HMC_CFG_GEAR_DOWN_EN (PRI_HMC_CFG_GEAR_DOWN_EN),
      .PRI_HMC_CFG_RLD3_MULTIBANK_MODE (PRI_HMC_CFG_RLD3_MULTIBANK_MODE),
      .PRI_HMC_CFG_PING_PONG_MODE (PRI_HMC_CFG_PING_PONG_MODE),
      .PRI_HMC_CFG_SLOT_ROTATE_EN (PRI_HMC_CFG_SLOT_ROTATE_EN),
      .PRI_HMC_CFG_SLOT_OFFSET (PRI_HMC_CFG_SLOT_OFFSET),
      .PRI_HMC_CFG_COL_CMD_SLOT (PRI_HMC_CFG_COL_CMD_SLOT),
      .PRI_HMC_CFG_ROW_CMD_SLOT (PRI_HMC_CFG_ROW_CMD_SLOT),
      .PRI_HMC_CFG_ENABLE_RC (PRI_HMC_CFG_ENABLE_RC),
      .PRI_HMC_CFG_CS_TO_CHIP_MAPPING (PRI_HMC_CFG_CS_TO_CHIP_MAPPING),
      .PRI_HMC_CFG_RB_RESERVED_ENTRY (PRI_HMC_CFG_RB_RESERVED_ENTRY),
      .PRI_HMC_CFG_WB_RESERVED_ENTRY (PRI_HMC_CFG_WB_RESERVED_ENTRY),
      .PRI_HMC_CFG_TCL (PRI_HMC_CFG_TCL),
      .PRI_HMC_CFG_POWER_SAVING_EXIT_CYC (PRI_HMC_CFG_POWER_SAVING_EXIT_CYC),
      .PRI_HMC_CFG_MEM_CLK_DISABLE_ENTRY_CYC (PRI_HMC_CFG_MEM_CLK_DISABLE_ENTRY_CYC),
      .PRI_HMC_CFG_WRITE_ODT_CHIP (PRI_HMC_CFG_WRITE_ODT_CHIP),
      .PRI_HMC_CFG_READ_ODT_CHIP (PRI_HMC_CFG_READ_ODT_CHIP),
      .PRI_HMC_CFG_WR_ODT_ON (PRI_HMC_CFG_WR_ODT_ON),
      .PRI_HMC_CFG_RD_ODT_ON (PRI_HMC_CFG_RD_ODT_ON),
      .PRI_HMC_CFG_WR_ODT_PERIOD (PRI_HMC_CFG_WR_ODT_PERIOD),
      .PRI_HMC_CFG_RD_ODT_PERIOD (PRI_HMC_CFG_RD_ODT_PERIOD),
      .PRI_HMC_CFG_RLD3_REFRESH_SEQ0 (PRI_HMC_CFG_RLD3_REFRESH_SEQ0),
      .PRI_HMC_CFG_RLD3_REFRESH_SEQ1 (PRI_HMC_CFG_RLD3_REFRESH_SEQ1),
      .PRI_HMC_CFG_RLD3_REFRESH_SEQ2 (PRI_HMC_CFG_RLD3_REFRESH_SEQ2),
      .PRI_HMC_CFG_RLD3_REFRESH_SEQ3 (PRI_HMC_CFG_RLD3_REFRESH_SEQ3),
      .PRI_HMC_CFG_SRF_ZQCAL_DISABLE (PRI_HMC_CFG_SRF_ZQCAL_DISABLE),
      .PRI_HMC_CFG_MPS_ZQCAL_DISABLE (PRI_HMC_CFG_MPS_ZQCAL_DISABLE),
      .PRI_HMC_CFG_MPS_DQSTRK_DISABLE (PRI_HMC_CFG_MPS_DQSTRK_DISABLE),
      .PRI_HMC_CFG_SHORT_DQSTRK_CTRL_EN (PRI_HMC_CFG_SHORT_DQSTRK_CTRL_EN),
      .PRI_HMC_CFG_PERIOD_DQSTRK_CTRL_EN (PRI_HMC_CFG_PERIOD_DQSTRK_CTRL_EN),
      .PRI_HMC_CFG_PERIOD_DQSTRK_INTERVAL (PRI_HMC_CFG_PERIOD_DQSTRK_INTERVAL),
      .PRI_HMC_CFG_DQSTRK_TO_VALID_LAST (PRI_HMC_CFG_DQSTRK_TO_VALID_LAST),
      .PRI_HMC_CFG_DQSTRK_TO_VALID (PRI_HMC_CFG_DQSTRK_TO_VALID),
      .PRI_HMC_CFG_RFSH_WARN_THRESHOLD (PRI_HMC_CFG_RFSH_WARN_THRESHOLD),
      .PRI_HMC_CFG_SB_CG_DISABLE (PRI_HMC_CFG_SB_CG_DISABLE),
      .PRI_HMC_CFG_USER_RFSH_EN (PRI_HMC_CFG_USER_RFSH_EN),
      .PRI_HMC_CFG_SRF_AUTOEXIT_EN (PRI_HMC_CFG_SRF_AUTOEXIT_EN),
      .PRI_HMC_CFG_SRF_ENTRY_EXIT_BLOCK (PRI_HMC_CFG_SRF_ENTRY_EXIT_BLOCK),
      .PRI_HMC_CFG_SB_DDR4_MR3 (PRI_HMC_CFG_SB_DDR4_MR3),
      .PRI_HMC_CFG_SB_DDR4_MR4 (PRI_HMC_CFG_SB_DDR4_MR4),
      .PRI_HMC_CFG_SB_DDR4_MR5 (PRI_HMC_CFG_SB_DDR4_MR5),
      .PRI_HMC_CFG_DDR4_MPS_ADDR_MIRROR (PRI_HMC_CFG_DDR4_MPS_ADDR_MIRROR),
      .PRI_HMC_CFG_MEM_IF_COLADDR_WIDTH (PRI_HMC_CFG_MEM_IF_COLADDR_WIDTH),
      .PRI_HMC_CFG_MEM_IF_ROWADDR_WIDTH (PRI_HMC_CFG_MEM_IF_ROWADDR_WIDTH),
      .PRI_HMC_CFG_MEM_IF_BANKADDR_WIDTH (PRI_HMC_CFG_MEM_IF_BANKADDR_WIDTH),
      .PRI_HMC_CFG_MEM_IF_BGADDR_WIDTH (PRI_HMC_CFG_MEM_IF_BGADDR_WIDTH),
      .PRI_HMC_CFG_LOCAL_IF_CS_WIDTH (PRI_HMC_CFG_LOCAL_IF_CS_WIDTH),
      .PRI_HMC_CFG_ADDR_ORDER (PRI_HMC_CFG_ADDR_ORDER),
      .PRI_HMC_CFG_ACT_TO_RDWR (PRI_HMC_CFG_ACT_TO_RDWR),
      .PRI_HMC_CFG_ACT_TO_PCH (PRI_HMC_CFG_ACT_TO_PCH),
      .PRI_HMC_CFG_ACT_TO_ACT (PRI_HMC_CFG_ACT_TO_ACT),
      .PRI_HMC_CFG_ACT_TO_ACT_DIFF_BANK (PRI_HMC_CFG_ACT_TO_ACT_DIFF_BANK),
      .PRI_HMC_CFG_ACT_TO_ACT_DIFF_BG (PRI_HMC_CFG_ACT_TO_ACT_DIFF_BG),
      .PRI_HMC_CFG_RD_TO_RD (PRI_HMC_CFG_RD_TO_RD),
      .PRI_HMC_CFG_RD_TO_RD_DIFF_CHIP (PRI_HMC_CFG_RD_TO_RD_DIFF_CHIP),
      .PRI_HMC_CFG_RD_TO_RD_DIFF_BG (PRI_HMC_CFG_RD_TO_RD_DIFF_BG),
      .PRI_HMC_CFG_RD_TO_WR (PRI_HMC_CFG_RD_TO_WR),
      .PRI_HMC_CFG_RD_TO_WR_DIFF_CHIP (PRI_HMC_CFG_RD_TO_WR_DIFF_CHIP),
      .PRI_HMC_CFG_RD_TO_WR_DIFF_BG (PRI_HMC_CFG_RD_TO_WR_DIFF_BG),
      .PRI_HMC_CFG_RD_TO_PCH (PRI_HMC_CFG_RD_TO_PCH),
      .PRI_HMC_CFG_RD_AP_TO_VALID (PRI_HMC_CFG_RD_AP_TO_VALID),
      .PRI_HMC_CFG_WR_TO_WR (PRI_HMC_CFG_WR_TO_WR),
      .PRI_HMC_CFG_WR_TO_WR_DIFF_CHIP (PRI_HMC_CFG_WR_TO_WR_DIFF_CHIP),
      .PRI_HMC_CFG_WR_TO_WR_DIFF_BG (PRI_HMC_CFG_WR_TO_WR_DIFF_BG),
      .PRI_HMC_CFG_WR_TO_RD (PRI_HMC_CFG_WR_TO_RD),
      .PRI_HMC_CFG_WR_TO_RD_DIFF_CHIP (PRI_HMC_CFG_WR_TO_RD_DIFF_CHIP),
      .PRI_HMC_CFG_WR_TO_RD_DIFF_BG (PRI_HMC_CFG_WR_TO_RD_DIFF_BG),
      .PRI_HMC_CFG_WR_TO_PCH (PRI_HMC_CFG_WR_TO_PCH),
      .PRI_HMC_CFG_WR_AP_TO_VALID (PRI_HMC_CFG_WR_AP_TO_VALID),
      .PRI_HMC_CFG_PCH_TO_VALID (PRI_HMC_CFG_PCH_TO_VALID),
      .PRI_HMC_CFG_PCH_ALL_TO_VALID (PRI_HMC_CFG_PCH_ALL_TO_VALID),
      .PRI_HMC_CFG_ARF_TO_VALID (PRI_HMC_CFG_ARF_TO_VALID),
      .PRI_HMC_CFG_PDN_TO_VALID (PRI_HMC_CFG_PDN_TO_VALID),
      .PRI_HMC_CFG_SRF_TO_VALID (PRI_HMC_CFG_SRF_TO_VALID),
      .PRI_HMC_CFG_SRF_TO_ZQ_CAL (PRI_HMC_CFG_SRF_TO_ZQ_CAL),
      .PRI_HMC_CFG_ARF_PERIOD (PRI_HMC_CFG_ARF_PERIOD),
      .PRI_HMC_CFG_PDN_PERIOD (PRI_HMC_CFG_PDN_PERIOD),
      .PRI_HMC_CFG_ZQCL_TO_VALID (PRI_HMC_CFG_ZQCL_TO_VALID),
      .PRI_HMC_CFG_ZQCS_TO_VALID (PRI_HMC_CFG_ZQCS_TO_VALID),
      .PRI_HMC_CFG_MRS_TO_VALID (PRI_HMC_CFG_MRS_TO_VALID),
      .PRI_HMC_CFG_MPS_TO_VALID (PRI_HMC_CFG_MPS_TO_VALID),
      .PRI_HMC_CFG_MRR_TO_VALID (PRI_HMC_CFG_MRR_TO_VALID),
      .PRI_HMC_CFG_MPR_TO_VALID (PRI_HMC_CFG_MPR_TO_VALID),
      .PRI_HMC_CFG_MPS_EXIT_CS_TO_CKE (PRI_HMC_CFG_MPS_EXIT_CS_TO_CKE),
      .PRI_HMC_CFG_MPS_EXIT_CKE_TO_CS (PRI_HMC_CFG_MPS_EXIT_CKE_TO_CS),
      .PRI_HMC_CFG_RLD3_MULTIBANK_REF_DELAY (PRI_HMC_CFG_RLD3_MULTIBANK_REF_DELAY),
      .PRI_HMC_CFG_MMR_CMD_TO_VALID (PRI_HMC_CFG_MMR_CMD_TO_VALID),
      .PRI_HMC_CFG_4_ACT_TO_ACT (PRI_HMC_CFG_4_ACT_TO_ACT),
      .PRI_HMC_CFG_16_ACT_TO_ACT (PRI_HMC_CFG_16_ACT_TO_ACT),
      .SEC_HMC_CFG_ENABLE_ECC (SEC_HMC_CFG_ENABLE_ECC),
      .SEC_HMC_CFG_REORDER_DATA (SEC_HMC_CFG_REORDER_DATA),
      .SEC_HMC_CFG_REORDER_READ (SEC_HMC_CFG_REORDER_READ),
      .SEC_HMC_CFG_REORDER_RDATA (SEC_HMC_CFG_REORDER_RDATA),
      .SEC_HMC_CFG_STARVE_LIMIT (SEC_HMC_CFG_STARVE_LIMIT),
      .SEC_HMC_CFG_DQS_TRACKING_EN (SEC_HMC_CFG_DQS_TRACKING_EN),
      .SEC_HMC_CFG_ARBITER_TYPE (SEC_HMC_CFG_ARBITER_TYPE),
      .SEC_HMC_CFG_OPEN_PAGE_EN (SEC_HMC_CFG_OPEN_PAGE_EN),
      .SEC_HMC_CFG_GEAR_DOWN_EN (SEC_HMC_CFG_GEAR_DOWN_EN),
      .SEC_HMC_CFG_RLD3_MULTIBANK_MODE (SEC_HMC_CFG_RLD3_MULTIBANK_MODE),
      .SEC_HMC_CFG_PING_PONG_MODE (SEC_HMC_CFG_PING_PONG_MODE),
      .SEC_HMC_CFG_SLOT_ROTATE_EN (SEC_HMC_CFG_SLOT_ROTATE_EN),
      .SEC_HMC_CFG_SLOT_OFFSET (SEC_HMC_CFG_SLOT_OFFSET),
      .SEC_HMC_CFG_COL_CMD_SLOT (SEC_HMC_CFG_COL_CMD_SLOT),
      .SEC_HMC_CFG_ROW_CMD_SLOT (SEC_HMC_CFG_ROW_CMD_SLOT),
      .SEC_HMC_CFG_ENABLE_RC (SEC_HMC_CFG_ENABLE_RC),
      .SEC_HMC_CFG_CS_TO_CHIP_MAPPING (SEC_HMC_CFG_CS_TO_CHIP_MAPPING),
      .SEC_HMC_CFG_RB_RESERVED_ENTRY (SEC_HMC_CFG_RB_RESERVED_ENTRY),
      .SEC_HMC_CFG_WB_RESERVED_ENTRY (SEC_HMC_CFG_WB_RESERVED_ENTRY),
      .SEC_HMC_CFG_TCL (SEC_HMC_CFG_TCL),
      .SEC_HMC_CFG_POWER_SAVING_EXIT_CYC (SEC_HMC_CFG_POWER_SAVING_EXIT_CYC),
      .SEC_HMC_CFG_MEM_CLK_DISABLE_ENTRY_CYC (SEC_HMC_CFG_MEM_CLK_DISABLE_ENTRY_CYC),
      .SEC_HMC_CFG_WRITE_ODT_CHIP (SEC_HMC_CFG_WRITE_ODT_CHIP),
      .SEC_HMC_CFG_READ_ODT_CHIP (SEC_HMC_CFG_READ_ODT_CHIP),
      .SEC_HMC_CFG_WR_ODT_ON (SEC_HMC_CFG_WR_ODT_ON),
      .SEC_HMC_CFG_RD_ODT_ON (SEC_HMC_CFG_RD_ODT_ON),
      .SEC_HMC_CFG_WR_ODT_PERIOD (SEC_HMC_CFG_WR_ODT_PERIOD),
      .SEC_HMC_CFG_RD_ODT_PERIOD (SEC_HMC_CFG_RD_ODT_PERIOD),
      .SEC_HMC_CFG_RLD3_REFRESH_SEQ0 (SEC_HMC_CFG_RLD3_REFRESH_SEQ0),
      .SEC_HMC_CFG_RLD3_REFRESH_SEQ1 (SEC_HMC_CFG_RLD3_REFRESH_SEQ1),
      .SEC_HMC_CFG_RLD3_REFRESH_SEQ2 (SEC_HMC_CFG_RLD3_REFRESH_SEQ2),
      .SEC_HMC_CFG_RLD3_REFRESH_SEQ3 (SEC_HMC_CFG_RLD3_REFRESH_SEQ3),
      .SEC_HMC_CFG_SRF_ZQCAL_DISABLE (SEC_HMC_CFG_SRF_ZQCAL_DISABLE),
      .SEC_HMC_CFG_MPS_ZQCAL_DISABLE (SEC_HMC_CFG_MPS_ZQCAL_DISABLE),
      .SEC_HMC_CFG_MPS_DQSTRK_DISABLE (SEC_HMC_CFG_MPS_DQSTRK_DISABLE),
      .SEC_HMC_CFG_SHORT_DQSTRK_CTRL_EN (SEC_HMC_CFG_SHORT_DQSTRK_CTRL_EN),
      .SEC_HMC_CFG_PERIOD_DQSTRK_CTRL_EN (SEC_HMC_CFG_PERIOD_DQSTRK_CTRL_EN),
      .SEC_HMC_CFG_PERIOD_DQSTRK_INTERVAL (SEC_HMC_CFG_PERIOD_DQSTRK_INTERVAL),
      .SEC_HMC_CFG_DQSTRK_TO_VALID_LAST (SEC_HMC_CFG_DQSTRK_TO_VALID_LAST),
      .SEC_HMC_CFG_DQSTRK_TO_VALID (SEC_HMC_CFG_DQSTRK_TO_VALID),
      .SEC_HMC_CFG_RFSH_WARN_THRESHOLD (SEC_HMC_CFG_RFSH_WARN_THRESHOLD),
      .SEC_HMC_CFG_SB_CG_DISABLE (SEC_HMC_CFG_SB_CG_DISABLE),
      .SEC_HMC_CFG_USER_RFSH_EN (SEC_HMC_CFG_USER_RFSH_EN),
      .SEC_HMC_CFG_SRF_AUTOEXIT_EN (SEC_HMC_CFG_SRF_AUTOEXIT_EN),
      .SEC_HMC_CFG_SRF_ENTRY_EXIT_BLOCK (SEC_HMC_CFG_SRF_ENTRY_EXIT_BLOCK),
      .SEC_HMC_CFG_SB_DDR4_MR3 (SEC_HMC_CFG_SB_DDR4_MR3),
      .SEC_HMC_CFG_SB_DDR4_MR4 (SEC_HMC_CFG_SB_DDR4_MR4),
      .SEC_HMC_CFG_SB_DDR4_MR5 (SEC_HMC_CFG_SB_DDR4_MR5),
      .SEC_HMC_CFG_DDR4_MPS_ADDR_MIRROR (SEC_HMC_CFG_DDR4_MPS_ADDR_MIRROR),
      .SEC_HMC_CFG_MEM_IF_COLADDR_WIDTH (SEC_HMC_CFG_MEM_IF_COLADDR_WIDTH),
      .SEC_HMC_CFG_MEM_IF_ROWADDR_WIDTH (SEC_HMC_CFG_MEM_IF_ROWADDR_WIDTH),
      .SEC_HMC_CFG_MEM_IF_BANKADDR_WIDTH (SEC_HMC_CFG_MEM_IF_BANKADDR_WIDTH),
      .SEC_HMC_CFG_MEM_IF_BGADDR_WIDTH (SEC_HMC_CFG_MEM_IF_BGADDR_WIDTH),
      .SEC_HMC_CFG_LOCAL_IF_CS_WIDTH (SEC_HMC_CFG_LOCAL_IF_CS_WIDTH),
      .SEC_HMC_CFG_ADDR_ORDER (SEC_HMC_CFG_ADDR_ORDER),
      .SEC_HMC_CFG_ACT_TO_RDWR (SEC_HMC_CFG_ACT_TO_RDWR),
      .SEC_HMC_CFG_ACT_TO_PCH (SEC_HMC_CFG_ACT_TO_PCH),
      .SEC_HMC_CFG_ACT_TO_ACT (SEC_HMC_CFG_ACT_TO_ACT),
      .SEC_HMC_CFG_ACT_TO_ACT_DIFF_BANK (SEC_HMC_CFG_ACT_TO_ACT_DIFF_BANK),
      .SEC_HMC_CFG_ACT_TO_ACT_DIFF_BG (SEC_HMC_CFG_ACT_TO_ACT_DIFF_BG),
      .SEC_HMC_CFG_RD_TO_RD (SEC_HMC_CFG_RD_TO_RD),
      .SEC_HMC_CFG_RD_TO_RD_DIFF_CHIP (SEC_HMC_CFG_RD_TO_RD_DIFF_CHIP),
      .SEC_HMC_CFG_RD_TO_RD_DIFF_BG (SEC_HMC_CFG_RD_TO_RD_DIFF_BG),
      .SEC_HMC_CFG_RD_TO_WR (SEC_HMC_CFG_RD_TO_WR),
      .SEC_HMC_CFG_RD_TO_WR_DIFF_CHIP (SEC_HMC_CFG_RD_TO_WR_DIFF_CHIP),
      .SEC_HMC_CFG_RD_TO_WR_DIFF_BG (SEC_HMC_CFG_RD_TO_WR_DIFF_BG),
      .SEC_HMC_CFG_RD_TO_PCH (SEC_HMC_CFG_RD_TO_PCH),
      .SEC_HMC_CFG_RD_AP_TO_VALID (SEC_HMC_CFG_RD_AP_TO_VALID),
      .SEC_HMC_CFG_WR_TO_WR (SEC_HMC_CFG_WR_TO_WR),
      .SEC_HMC_CFG_WR_TO_WR_DIFF_CHIP (SEC_HMC_CFG_WR_TO_WR_DIFF_CHIP),
      .SEC_HMC_CFG_WR_TO_WR_DIFF_BG (SEC_HMC_CFG_WR_TO_WR_DIFF_BG),
      .SEC_HMC_CFG_WR_TO_RD (SEC_HMC_CFG_WR_TO_RD),
      .SEC_HMC_CFG_WR_TO_RD_DIFF_CHIP (SEC_HMC_CFG_WR_TO_RD_DIFF_CHIP),
      .SEC_HMC_CFG_WR_TO_RD_DIFF_BG (SEC_HMC_CFG_WR_TO_RD_DIFF_BG),
      .SEC_HMC_CFG_WR_TO_PCH (SEC_HMC_CFG_WR_TO_PCH),
      .SEC_HMC_CFG_WR_AP_TO_VALID (SEC_HMC_CFG_WR_AP_TO_VALID),
      .SEC_HMC_CFG_PCH_TO_VALID (SEC_HMC_CFG_PCH_TO_VALID),
      .SEC_HMC_CFG_PCH_ALL_TO_VALID (SEC_HMC_CFG_PCH_ALL_TO_VALID),
      .SEC_HMC_CFG_ARF_TO_VALID (SEC_HMC_CFG_ARF_TO_VALID),
      .SEC_HMC_CFG_PDN_TO_VALID (SEC_HMC_CFG_PDN_TO_VALID),
      .SEC_HMC_CFG_SRF_TO_VALID (SEC_HMC_CFG_SRF_TO_VALID),
      .SEC_HMC_CFG_SRF_TO_ZQ_CAL (SEC_HMC_CFG_SRF_TO_ZQ_CAL),
      .SEC_HMC_CFG_ARF_PERIOD (SEC_HMC_CFG_ARF_PERIOD),
      .SEC_HMC_CFG_PDN_PERIOD (SEC_HMC_CFG_PDN_PERIOD),
      .SEC_HMC_CFG_ZQCL_TO_VALID (SEC_HMC_CFG_ZQCL_TO_VALID),
      .SEC_HMC_CFG_ZQCS_TO_VALID (SEC_HMC_CFG_ZQCS_TO_VALID),
      .SEC_HMC_CFG_MRS_TO_VALID (SEC_HMC_CFG_MRS_TO_VALID),
      .SEC_HMC_CFG_MPS_TO_VALID (SEC_HMC_CFG_MPS_TO_VALID),
      .SEC_HMC_CFG_MRR_TO_VALID (SEC_HMC_CFG_MRR_TO_VALID),
      .SEC_HMC_CFG_MPR_TO_VALID (SEC_HMC_CFG_MPR_TO_VALID),
      .SEC_HMC_CFG_MPS_EXIT_CS_TO_CKE (SEC_HMC_CFG_MPS_EXIT_CS_TO_CKE),
      .SEC_HMC_CFG_MPS_EXIT_CKE_TO_CS (SEC_HMC_CFG_MPS_EXIT_CKE_TO_CS),
      .SEC_HMC_CFG_RLD3_MULTIBANK_REF_DELAY (SEC_HMC_CFG_RLD3_MULTIBANK_REF_DELAY),
      .SEC_HMC_CFG_MMR_CMD_TO_VALID (SEC_HMC_CFG_MMR_CMD_TO_VALID),
      .SEC_HMC_CFG_4_ACT_TO_ACT (SEC_HMC_CFG_4_ACT_TO_ACT),
      .SEC_HMC_CFG_16_ACT_TO_ACT (SEC_HMC_CFG_16_ACT_TO_ACT),
      .PINS_PER_LANE (PINS_PER_LANE),
      .LANES_PER_TILE (LANES_PER_TILE),
      .OCT_CONTROL_WIDTH (OCT_CONTROL_WIDTH),
      .PORT_MEM_CK_WIDTH (PORT_MEM_CK_WIDTH),
      .PORT_MEM_CK_PINLOC_0 (PORT_MEM_CK_PINLOC_0),
      .PORT_MEM_CK_PINLOC_1 (PORT_MEM_CK_PINLOC_1),
      .PORT_MEM_CK_PINLOC_2 (PORT_MEM_CK_PINLOC_2),
      .PORT_MEM_CK_PINLOC_3 (PORT_MEM_CK_PINLOC_3),
      .PORT_MEM_CK_PINLOC_4 (PORT_MEM_CK_PINLOC_4),
      .PORT_MEM_CK_PINLOC_5 (PORT_MEM_CK_PINLOC_5),
      .PORT_MEM_CK_PINLOC_AUTOGEN_WCNT (PORT_MEM_CK_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CK_N_WIDTH (PORT_MEM_CK_N_WIDTH),
      .PORT_MEM_CK_N_PINLOC_0 (PORT_MEM_CK_N_PINLOC_0),
      .PORT_MEM_CK_N_PINLOC_1 (PORT_MEM_CK_N_PINLOC_1),
      .PORT_MEM_CK_N_PINLOC_2 (PORT_MEM_CK_N_PINLOC_2),
      .PORT_MEM_CK_N_PINLOC_3 (PORT_MEM_CK_N_PINLOC_3),
      .PORT_MEM_CK_N_PINLOC_4 (PORT_MEM_CK_N_PINLOC_4),
      .PORT_MEM_CK_N_PINLOC_5 (PORT_MEM_CK_N_PINLOC_5),
      .PORT_MEM_CK_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_CK_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DK_WIDTH (PORT_MEM_DK_WIDTH),
      .PORT_MEM_DK_PINLOC_0 (PORT_MEM_DK_PINLOC_0),
      .PORT_MEM_DK_PINLOC_1 (PORT_MEM_DK_PINLOC_1),
      .PORT_MEM_DK_PINLOC_2 (PORT_MEM_DK_PINLOC_2),
      .PORT_MEM_DK_PINLOC_3 (PORT_MEM_DK_PINLOC_3),
      .PORT_MEM_DK_PINLOC_4 (PORT_MEM_DK_PINLOC_4),
      .PORT_MEM_DK_PINLOC_5 (PORT_MEM_DK_PINLOC_5),
      .PORT_MEM_DK_PINLOC_AUTOGEN_WCNT (PORT_MEM_DK_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DK_N_WIDTH (PORT_MEM_DK_N_WIDTH),
      .PORT_MEM_DK_N_PINLOC_0 (PORT_MEM_DK_N_PINLOC_0),
      .PORT_MEM_DK_N_PINLOC_1 (PORT_MEM_DK_N_PINLOC_1),
      .PORT_MEM_DK_N_PINLOC_2 (PORT_MEM_DK_N_PINLOC_2),
      .PORT_MEM_DK_N_PINLOC_3 (PORT_MEM_DK_N_PINLOC_3),
      .PORT_MEM_DK_N_PINLOC_4 (PORT_MEM_DK_N_PINLOC_4),
      .PORT_MEM_DK_N_PINLOC_5 (PORT_MEM_DK_N_PINLOC_5),
      .PORT_MEM_DK_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_DK_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DKA_WIDTH (PORT_MEM_DKA_WIDTH),
      .PORT_MEM_DKA_PINLOC_0 (PORT_MEM_DKA_PINLOC_0),
      .PORT_MEM_DKA_PINLOC_1 (PORT_MEM_DKA_PINLOC_1),
      .PORT_MEM_DKA_PINLOC_2 (PORT_MEM_DKA_PINLOC_2),
      .PORT_MEM_DKA_PINLOC_3 (PORT_MEM_DKA_PINLOC_3),
      .PORT_MEM_DKA_PINLOC_4 (PORT_MEM_DKA_PINLOC_4),
      .PORT_MEM_DKA_PINLOC_5 (PORT_MEM_DKA_PINLOC_5),
      .PORT_MEM_DKA_PINLOC_AUTOGEN_WCNT (PORT_MEM_DKA_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DKA_N_WIDTH (PORT_MEM_DKA_N_WIDTH),
      .PORT_MEM_DKA_N_PINLOC_0 (PORT_MEM_DKA_N_PINLOC_0),
      .PORT_MEM_DKA_N_PINLOC_1 (PORT_MEM_DKA_N_PINLOC_1),
      .PORT_MEM_DKA_N_PINLOC_2 (PORT_MEM_DKA_N_PINLOC_2),
      .PORT_MEM_DKA_N_PINLOC_3 (PORT_MEM_DKA_N_PINLOC_3),
      .PORT_MEM_DKA_N_PINLOC_4 (PORT_MEM_DKA_N_PINLOC_4),
      .PORT_MEM_DKA_N_PINLOC_5 (PORT_MEM_DKA_N_PINLOC_5),
      .PORT_MEM_DKA_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_DKA_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DKB_WIDTH (PORT_MEM_DKB_WIDTH),
      .PORT_MEM_DKB_PINLOC_0 (PORT_MEM_DKB_PINLOC_0),
      .PORT_MEM_DKB_PINLOC_1 (PORT_MEM_DKB_PINLOC_1),
      .PORT_MEM_DKB_PINLOC_2 (PORT_MEM_DKB_PINLOC_2),
      .PORT_MEM_DKB_PINLOC_3 (PORT_MEM_DKB_PINLOC_3),
      .PORT_MEM_DKB_PINLOC_4 (PORT_MEM_DKB_PINLOC_4),
      .PORT_MEM_DKB_PINLOC_5 (PORT_MEM_DKB_PINLOC_5),
      .PORT_MEM_DKB_PINLOC_AUTOGEN_WCNT (PORT_MEM_DKB_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DKB_N_WIDTH (PORT_MEM_DKB_N_WIDTH),
      .PORT_MEM_DKB_N_PINLOC_0 (PORT_MEM_DKB_N_PINLOC_0),
      .PORT_MEM_DKB_N_PINLOC_1 (PORT_MEM_DKB_N_PINLOC_1),
      .PORT_MEM_DKB_N_PINLOC_2 (PORT_MEM_DKB_N_PINLOC_2),
      .PORT_MEM_DKB_N_PINLOC_3 (PORT_MEM_DKB_N_PINLOC_3),
      .PORT_MEM_DKB_N_PINLOC_4 (PORT_MEM_DKB_N_PINLOC_4),
      .PORT_MEM_DKB_N_PINLOC_5 (PORT_MEM_DKB_N_PINLOC_5),
      .PORT_MEM_DKB_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_DKB_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_K_WIDTH (PORT_MEM_K_WIDTH),
      .PORT_MEM_K_PINLOC_0 (PORT_MEM_K_PINLOC_0),
      .PORT_MEM_K_PINLOC_1 (PORT_MEM_K_PINLOC_1),
      .PORT_MEM_K_PINLOC_2 (PORT_MEM_K_PINLOC_2),
      .PORT_MEM_K_PINLOC_3 (PORT_MEM_K_PINLOC_3),
      .PORT_MEM_K_PINLOC_4 (PORT_MEM_K_PINLOC_4),
      .PORT_MEM_K_PINLOC_5 (PORT_MEM_K_PINLOC_5),
      .PORT_MEM_K_PINLOC_AUTOGEN_WCNT (PORT_MEM_K_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_K_N_WIDTH (PORT_MEM_K_N_WIDTH),
      .PORT_MEM_K_N_PINLOC_0 (PORT_MEM_K_N_PINLOC_0),
      .PORT_MEM_K_N_PINLOC_1 (PORT_MEM_K_N_PINLOC_1),
      .PORT_MEM_K_N_PINLOC_2 (PORT_MEM_K_N_PINLOC_2),
      .PORT_MEM_K_N_PINLOC_3 (PORT_MEM_K_N_PINLOC_3),
      .PORT_MEM_K_N_PINLOC_4 (PORT_MEM_K_N_PINLOC_4),
      .PORT_MEM_K_N_PINLOC_5 (PORT_MEM_K_N_PINLOC_5),
      .PORT_MEM_K_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_K_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_A_WIDTH (PORT_MEM_A_WIDTH),
      .PORT_MEM_A_PINLOC_0 (PORT_MEM_A_PINLOC_0),
      .PORT_MEM_A_PINLOC_1 (PORT_MEM_A_PINLOC_1),
      .PORT_MEM_A_PINLOC_2 (PORT_MEM_A_PINLOC_2),
      .PORT_MEM_A_PINLOC_3 (PORT_MEM_A_PINLOC_3),
      .PORT_MEM_A_PINLOC_4 (PORT_MEM_A_PINLOC_4),
      .PORT_MEM_A_PINLOC_5 (PORT_MEM_A_PINLOC_5),
      .PORT_MEM_A_PINLOC_6 (PORT_MEM_A_PINLOC_6),
      .PORT_MEM_A_PINLOC_7 (PORT_MEM_A_PINLOC_7),
      .PORT_MEM_A_PINLOC_8 (PORT_MEM_A_PINLOC_8),
      .PORT_MEM_A_PINLOC_9 (PORT_MEM_A_PINLOC_9),
      .PORT_MEM_A_PINLOC_10 (PORT_MEM_A_PINLOC_10),
      .PORT_MEM_A_PINLOC_11 (PORT_MEM_A_PINLOC_11),
      .PORT_MEM_A_PINLOC_12 (PORT_MEM_A_PINLOC_12),
      .PORT_MEM_A_PINLOC_13 (PORT_MEM_A_PINLOC_13),
      .PORT_MEM_A_PINLOC_14 (PORT_MEM_A_PINLOC_14),
      .PORT_MEM_A_PINLOC_15 (PORT_MEM_A_PINLOC_15),
      .PORT_MEM_A_PINLOC_16 (PORT_MEM_A_PINLOC_16),
      .PORT_MEM_A_PINLOC_AUTOGEN_WCNT (PORT_MEM_A_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_BA_WIDTH (PORT_MEM_BA_WIDTH),
      .PORT_MEM_BA_PINLOC_0 (PORT_MEM_BA_PINLOC_0),
      .PORT_MEM_BA_PINLOC_1 (PORT_MEM_BA_PINLOC_1),
      .PORT_MEM_BA_PINLOC_2 (PORT_MEM_BA_PINLOC_2),
      .PORT_MEM_BA_PINLOC_3 (PORT_MEM_BA_PINLOC_3),
      .PORT_MEM_BA_PINLOC_4 (PORT_MEM_BA_PINLOC_4),
      .PORT_MEM_BA_PINLOC_5 (PORT_MEM_BA_PINLOC_5),
      .PORT_MEM_BA_PINLOC_AUTOGEN_WCNT (PORT_MEM_BA_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_BG_WIDTH (PORT_MEM_BG_WIDTH),
      .PORT_MEM_BG_PINLOC_0 (PORT_MEM_BG_PINLOC_0),
      .PORT_MEM_BG_PINLOC_1 (PORT_MEM_BG_PINLOC_1),
      .PORT_MEM_BG_PINLOC_2 (PORT_MEM_BG_PINLOC_2),
      .PORT_MEM_BG_PINLOC_3 (PORT_MEM_BG_PINLOC_3),
      .PORT_MEM_BG_PINLOC_4 (PORT_MEM_BG_PINLOC_4),
      .PORT_MEM_BG_PINLOC_5 (PORT_MEM_BG_PINLOC_5),
      .PORT_MEM_BG_PINLOC_AUTOGEN_WCNT (PORT_MEM_BG_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_C_WIDTH (PORT_MEM_C_WIDTH),
      .PORT_MEM_C_PINLOC_0 (PORT_MEM_C_PINLOC_0),
      .PORT_MEM_C_PINLOC_1 (PORT_MEM_C_PINLOC_1),
      .PORT_MEM_C_PINLOC_2 (PORT_MEM_C_PINLOC_2),
      .PORT_MEM_C_PINLOC_3 (PORT_MEM_C_PINLOC_3),
      .PORT_MEM_C_PINLOC_4 (PORT_MEM_C_PINLOC_4),
      .PORT_MEM_C_PINLOC_5 (PORT_MEM_C_PINLOC_5),
      .PORT_MEM_C_PINLOC_AUTOGEN_WCNT (PORT_MEM_C_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CKE_WIDTH (PORT_MEM_CKE_WIDTH),
      .PORT_MEM_CKE_PINLOC_0 (PORT_MEM_CKE_PINLOC_0),
      .PORT_MEM_CKE_PINLOC_1 (PORT_MEM_CKE_PINLOC_1),
      .PORT_MEM_CKE_PINLOC_2 (PORT_MEM_CKE_PINLOC_2),
      .PORT_MEM_CKE_PINLOC_3 (PORT_MEM_CKE_PINLOC_3),
      .PORT_MEM_CKE_PINLOC_4 (PORT_MEM_CKE_PINLOC_4),
      .PORT_MEM_CKE_PINLOC_5 (PORT_MEM_CKE_PINLOC_5),
      .PORT_MEM_CKE_PINLOC_AUTOGEN_WCNT (PORT_MEM_CKE_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CS_N_WIDTH (PORT_MEM_CS_N_WIDTH),
      .PORT_MEM_CS_N_PINLOC_0 (PORT_MEM_CS_N_PINLOC_0),
      .PORT_MEM_CS_N_PINLOC_1 (PORT_MEM_CS_N_PINLOC_1),
      .PORT_MEM_CS_N_PINLOC_2 (PORT_MEM_CS_N_PINLOC_2),
      .PORT_MEM_CS_N_PINLOC_3 (PORT_MEM_CS_N_PINLOC_3),
      .PORT_MEM_CS_N_PINLOC_4 (PORT_MEM_CS_N_PINLOC_4),
      .PORT_MEM_CS_N_PINLOC_5 (PORT_MEM_CS_N_PINLOC_5),
      .PORT_MEM_CS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_CS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_RM_WIDTH (PORT_MEM_RM_WIDTH),
      .PORT_MEM_RM_PINLOC_0 (PORT_MEM_RM_PINLOC_0),
      .PORT_MEM_RM_PINLOC_1 (PORT_MEM_RM_PINLOC_1),
      .PORT_MEM_RM_PINLOC_2 (PORT_MEM_RM_PINLOC_2),
      .PORT_MEM_RM_PINLOC_3 (PORT_MEM_RM_PINLOC_3),
      .PORT_MEM_RM_PINLOC_4 (PORT_MEM_RM_PINLOC_4),
      .PORT_MEM_RM_PINLOC_5 (PORT_MEM_RM_PINLOC_5),
      .PORT_MEM_RM_PINLOC_AUTOGEN_WCNT (PORT_MEM_RM_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_ODT_WIDTH (PORT_MEM_ODT_WIDTH),
      .PORT_MEM_ODT_PINLOC_0 (PORT_MEM_ODT_PINLOC_0),
      .PORT_MEM_ODT_PINLOC_1 (PORT_MEM_ODT_PINLOC_1),
      .PORT_MEM_ODT_PINLOC_2 (PORT_MEM_ODT_PINLOC_2),
      .PORT_MEM_ODT_PINLOC_3 (PORT_MEM_ODT_PINLOC_3),
      .PORT_MEM_ODT_PINLOC_4 (PORT_MEM_ODT_PINLOC_4),
      .PORT_MEM_ODT_PINLOC_5 (PORT_MEM_ODT_PINLOC_5),
      .PORT_MEM_ODT_PINLOC_AUTOGEN_WCNT (PORT_MEM_ODT_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_RAS_N_WIDTH (PORT_MEM_RAS_N_WIDTH),
      .PORT_MEM_RAS_N_PINLOC_0 (PORT_MEM_RAS_N_PINLOC_0),
      .PORT_MEM_RAS_N_PINLOC_1 (PORT_MEM_RAS_N_PINLOC_1),
      .PORT_MEM_RAS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_RAS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CAS_N_WIDTH (PORT_MEM_CAS_N_WIDTH),
      .PORT_MEM_CAS_N_PINLOC_0 (PORT_MEM_CAS_N_PINLOC_0),
      .PORT_MEM_CAS_N_PINLOC_1 (PORT_MEM_CAS_N_PINLOC_1),
      .PORT_MEM_CAS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_CAS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_WE_N_WIDTH (PORT_MEM_WE_N_WIDTH),
      .PORT_MEM_WE_N_PINLOC_0 (PORT_MEM_WE_N_PINLOC_0),
      .PORT_MEM_WE_N_PINLOC_1 (PORT_MEM_WE_N_PINLOC_1),
      .PORT_MEM_WE_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_WE_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_RESET_N_WIDTH (PORT_MEM_RESET_N_WIDTH),
      .PORT_MEM_RESET_N_PINLOC_0 (PORT_MEM_RESET_N_PINLOC_0),
      .PORT_MEM_RESET_N_PINLOC_1 (PORT_MEM_RESET_N_PINLOC_1),
      .PORT_MEM_RESET_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_RESET_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_ACT_N_WIDTH (PORT_MEM_ACT_N_WIDTH),
      .PORT_MEM_ACT_N_PINLOC_0 (PORT_MEM_ACT_N_PINLOC_0),
      .PORT_MEM_ACT_N_PINLOC_1 (PORT_MEM_ACT_N_PINLOC_1),
      .PORT_MEM_ACT_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_ACT_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_PAR_WIDTH (PORT_MEM_PAR_WIDTH),
      .PORT_MEM_PAR_PINLOC_0 (PORT_MEM_PAR_PINLOC_0),
      .PORT_MEM_PAR_PINLOC_1 (PORT_MEM_PAR_PINLOC_1),
      .PORT_MEM_PAR_PINLOC_AUTOGEN_WCNT (PORT_MEM_PAR_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CA_WIDTH (PORT_MEM_CA_WIDTH),
      .PORT_MEM_CA_PINLOC_0 (PORT_MEM_CA_PINLOC_0),
      .PORT_MEM_CA_PINLOC_1 (PORT_MEM_CA_PINLOC_1),
      .PORT_MEM_CA_PINLOC_2 (PORT_MEM_CA_PINLOC_2),
      .PORT_MEM_CA_PINLOC_3 (PORT_MEM_CA_PINLOC_3),
      .PORT_MEM_CA_PINLOC_4 (PORT_MEM_CA_PINLOC_4),
      .PORT_MEM_CA_PINLOC_5 (PORT_MEM_CA_PINLOC_5),
      .PORT_MEM_CA_PINLOC_6 (PORT_MEM_CA_PINLOC_6),
      .PORT_MEM_CA_PINLOC_7 (PORT_MEM_CA_PINLOC_7),
      .PORT_MEM_CA_PINLOC_8 (PORT_MEM_CA_PINLOC_8),
      .PORT_MEM_CA_PINLOC_9 (PORT_MEM_CA_PINLOC_9),
      .PORT_MEM_CA_PINLOC_10 (PORT_MEM_CA_PINLOC_10),
      .PORT_MEM_CA_PINLOC_11 (PORT_MEM_CA_PINLOC_11),
      .PORT_MEM_CA_PINLOC_12 (PORT_MEM_CA_PINLOC_12),
      .PORT_MEM_CA_PINLOC_13 (PORT_MEM_CA_PINLOC_13),
      .PORT_MEM_CA_PINLOC_14 (PORT_MEM_CA_PINLOC_14),
      .PORT_MEM_CA_PINLOC_15 (PORT_MEM_CA_PINLOC_15),
      .PORT_MEM_CA_PINLOC_16 (PORT_MEM_CA_PINLOC_16),
      .PORT_MEM_CA_PINLOC_AUTOGEN_WCNT (PORT_MEM_CA_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_REF_N_WIDTH (PORT_MEM_REF_N_WIDTH),
      .PORT_MEM_REF_N_PINLOC_0 (PORT_MEM_REF_N_PINLOC_0),
      .PORT_MEM_REF_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_REF_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_WPS_N_WIDTH (PORT_MEM_WPS_N_WIDTH),
      .PORT_MEM_WPS_N_PINLOC_0 (PORT_MEM_WPS_N_PINLOC_0),
      .PORT_MEM_WPS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_WPS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_RPS_N_WIDTH (PORT_MEM_RPS_N_WIDTH),
      .PORT_MEM_RPS_N_PINLOC_0 (PORT_MEM_RPS_N_PINLOC_0),
      .PORT_MEM_RPS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_RPS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DOFF_N_WIDTH (PORT_MEM_DOFF_N_WIDTH),
      .PORT_MEM_DOFF_N_PINLOC_0 (PORT_MEM_DOFF_N_PINLOC_0),
      .PORT_MEM_DOFF_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_DOFF_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_LDA_N_WIDTH (PORT_MEM_LDA_N_WIDTH),
      .PORT_MEM_LDA_N_PINLOC_0 (PORT_MEM_LDA_N_PINLOC_0),
      .PORT_MEM_LDA_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_LDA_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_LDB_N_WIDTH (PORT_MEM_LDB_N_WIDTH),
      .PORT_MEM_LDB_N_PINLOC_0 (PORT_MEM_LDB_N_PINLOC_0),
      .PORT_MEM_LDB_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_LDB_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_RWA_N_WIDTH (PORT_MEM_RWA_N_WIDTH),
      .PORT_MEM_RWA_N_PINLOC_0 (PORT_MEM_RWA_N_PINLOC_0),
      .PORT_MEM_RWA_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_RWA_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_RWB_N_WIDTH (PORT_MEM_RWB_N_WIDTH),
      .PORT_MEM_RWB_N_PINLOC_0 (PORT_MEM_RWB_N_PINLOC_0),
      .PORT_MEM_RWB_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_RWB_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_LBK0_N_WIDTH (PORT_MEM_LBK0_N_WIDTH),
      .PORT_MEM_LBK0_N_PINLOC_0 (PORT_MEM_LBK0_N_PINLOC_0),
      .PORT_MEM_LBK0_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_LBK0_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_LBK1_N_WIDTH (PORT_MEM_LBK1_N_WIDTH),
      .PORT_MEM_LBK1_N_PINLOC_0 (PORT_MEM_LBK1_N_PINLOC_0),
      .PORT_MEM_LBK1_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_LBK1_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CFG_N_WIDTH (PORT_MEM_CFG_N_WIDTH),
      .PORT_MEM_CFG_N_PINLOC_0 (PORT_MEM_CFG_N_PINLOC_0),
      .PORT_MEM_CFG_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_CFG_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_AP_WIDTH (PORT_MEM_AP_WIDTH),
      .PORT_MEM_AP_PINLOC_0 (PORT_MEM_AP_PINLOC_0),
      .PORT_MEM_AP_PINLOC_AUTOGEN_WCNT (PORT_MEM_AP_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_AINV_WIDTH (PORT_MEM_AINV_WIDTH),
      .PORT_MEM_AINV_PINLOC_0 (PORT_MEM_AINV_PINLOC_0),
      .PORT_MEM_AINV_PINLOC_AUTOGEN_WCNT (PORT_MEM_AINV_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DM_WIDTH (PORT_MEM_DM_WIDTH),
      .PORT_MEM_DM_PINLOC_0 (PORT_MEM_DM_PINLOC_0),
      .PORT_MEM_DM_PINLOC_1 (PORT_MEM_DM_PINLOC_1),
      .PORT_MEM_DM_PINLOC_2 (PORT_MEM_DM_PINLOC_2),
      .PORT_MEM_DM_PINLOC_3 (PORT_MEM_DM_PINLOC_3),
      .PORT_MEM_DM_PINLOC_4 (PORT_MEM_DM_PINLOC_4),
      .PORT_MEM_DM_PINLOC_5 (PORT_MEM_DM_PINLOC_5),
      .PORT_MEM_DM_PINLOC_6 (PORT_MEM_DM_PINLOC_6),
      .PORT_MEM_DM_PINLOC_7 (PORT_MEM_DM_PINLOC_7),
      .PORT_MEM_DM_PINLOC_8 (PORT_MEM_DM_PINLOC_8),
      .PORT_MEM_DM_PINLOC_9 (PORT_MEM_DM_PINLOC_9),
      .PORT_MEM_DM_PINLOC_10 (PORT_MEM_DM_PINLOC_10),
      .PORT_MEM_DM_PINLOC_11 (PORT_MEM_DM_PINLOC_11),
      .PORT_MEM_DM_PINLOC_12 (PORT_MEM_DM_PINLOC_12),
      .PORT_MEM_DM_PINLOC_AUTOGEN_WCNT (PORT_MEM_DM_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_BWS_N_WIDTH (PORT_MEM_BWS_N_WIDTH),
      .PORT_MEM_BWS_N_PINLOC_0 (PORT_MEM_BWS_N_PINLOC_0),
      .PORT_MEM_BWS_N_PINLOC_1 (PORT_MEM_BWS_N_PINLOC_1),
      .PORT_MEM_BWS_N_PINLOC_2 (PORT_MEM_BWS_N_PINLOC_2),
      .PORT_MEM_BWS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_BWS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_D_WIDTH (PORT_MEM_D_WIDTH),
      .PORT_MEM_D_PINLOC_0 (PORT_MEM_D_PINLOC_0),
      .PORT_MEM_D_PINLOC_1 (PORT_MEM_D_PINLOC_1),
      .PORT_MEM_D_PINLOC_2 (PORT_MEM_D_PINLOC_2),
      .PORT_MEM_D_PINLOC_3 (PORT_MEM_D_PINLOC_3),
      .PORT_MEM_D_PINLOC_4 (PORT_MEM_D_PINLOC_4),
      .PORT_MEM_D_PINLOC_5 (PORT_MEM_D_PINLOC_5),
      .PORT_MEM_D_PINLOC_6 (PORT_MEM_D_PINLOC_6),
      .PORT_MEM_D_PINLOC_7 (PORT_MEM_D_PINLOC_7),
      .PORT_MEM_D_PINLOC_8 (PORT_MEM_D_PINLOC_8),
      .PORT_MEM_D_PINLOC_9 (PORT_MEM_D_PINLOC_9),
      .PORT_MEM_D_PINLOC_10 (PORT_MEM_D_PINLOC_10),
      .PORT_MEM_D_PINLOC_11 (PORT_MEM_D_PINLOC_11),
      .PORT_MEM_D_PINLOC_12 (PORT_MEM_D_PINLOC_12),
      .PORT_MEM_D_PINLOC_13 (PORT_MEM_D_PINLOC_13),
      .PORT_MEM_D_PINLOC_14 (PORT_MEM_D_PINLOC_14),
      .PORT_MEM_D_PINLOC_15 (PORT_MEM_D_PINLOC_15),
      .PORT_MEM_D_PINLOC_16 (PORT_MEM_D_PINLOC_16),
      .PORT_MEM_D_PINLOC_17 (PORT_MEM_D_PINLOC_17),
      .PORT_MEM_D_PINLOC_18 (PORT_MEM_D_PINLOC_18),
      .PORT_MEM_D_PINLOC_19 (PORT_MEM_D_PINLOC_19),
      .PORT_MEM_D_PINLOC_20 (PORT_MEM_D_PINLOC_20),
      .PORT_MEM_D_PINLOC_21 (PORT_MEM_D_PINLOC_21),
      .PORT_MEM_D_PINLOC_22 (PORT_MEM_D_PINLOC_22),
      .PORT_MEM_D_PINLOC_23 (PORT_MEM_D_PINLOC_23),
      .PORT_MEM_D_PINLOC_24 (PORT_MEM_D_PINLOC_24),
      .PORT_MEM_D_PINLOC_25 (PORT_MEM_D_PINLOC_25),
      .PORT_MEM_D_PINLOC_26 (PORT_MEM_D_PINLOC_26),
      .PORT_MEM_D_PINLOC_27 (PORT_MEM_D_PINLOC_27),
      .PORT_MEM_D_PINLOC_28 (PORT_MEM_D_PINLOC_28),
      .PORT_MEM_D_PINLOC_29 (PORT_MEM_D_PINLOC_29),
      .PORT_MEM_D_PINLOC_30 (PORT_MEM_D_PINLOC_30),
      .PORT_MEM_D_PINLOC_31 (PORT_MEM_D_PINLOC_31),
      .PORT_MEM_D_PINLOC_32 (PORT_MEM_D_PINLOC_32),
      .PORT_MEM_D_PINLOC_33 (PORT_MEM_D_PINLOC_33),
      .PORT_MEM_D_PINLOC_34 (PORT_MEM_D_PINLOC_34),
      .PORT_MEM_D_PINLOC_35 (PORT_MEM_D_PINLOC_35),
      .PORT_MEM_D_PINLOC_36 (PORT_MEM_D_PINLOC_36),
      .PORT_MEM_D_PINLOC_37 (PORT_MEM_D_PINLOC_37),
      .PORT_MEM_D_PINLOC_38 (PORT_MEM_D_PINLOC_38),
      .PORT_MEM_D_PINLOC_39 (PORT_MEM_D_PINLOC_39),
      .PORT_MEM_D_PINLOC_40 (PORT_MEM_D_PINLOC_40),
      .PORT_MEM_D_PINLOC_41 (PORT_MEM_D_PINLOC_41),
      .PORT_MEM_D_PINLOC_42 (PORT_MEM_D_PINLOC_42),
      .PORT_MEM_D_PINLOC_43 (PORT_MEM_D_PINLOC_43),
      .PORT_MEM_D_PINLOC_44 (PORT_MEM_D_PINLOC_44),
      .PORT_MEM_D_PINLOC_45 (PORT_MEM_D_PINLOC_45),
      .PORT_MEM_D_PINLOC_46 (PORT_MEM_D_PINLOC_46),
      .PORT_MEM_D_PINLOC_47 (PORT_MEM_D_PINLOC_47),
      .PORT_MEM_D_PINLOC_48 (PORT_MEM_D_PINLOC_48),
      .PORT_MEM_D_PINLOC_AUTOGEN_WCNT (PORT_MEM_D_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DQ_WIDTH (PORT_MEM_DQ_WIDTH),
      .PORT_MEM_DQ_PINLOC_0 (PORT_MEM_DQ_PINLOC_0),
      .PORT_MEM_DQ_PINLOC_1 (PORT_MEM_DQ_PINLOC_1),
      .PORT_MEM_DQ_PINLOC_2 (PORT_MEM_DQ_PINLOC_2),
      .PORT_MEM_DQ_PINLOC_3 (PORT_MEM_DQ_PINLOC_3),
      .PORT_MEM_DQ_PINLOC_4 (PORT_MEM_DQ_PINLOC_4),
      .PORT_MEM_DQ_PINLOC_5 (PORT_MEM_DQ_PINLOC_5),
      .PORT_MEM_DQ_PINLOC_6 (PORT_MEM_DQ_PINLOC_6),
      .PORT_MEM_DQ_PINLOC_7 (PORT_MEM_DQ_PINLOC_7),
      .PORT_MEM_DQ_PINLOC_8 (PORT_MEM_DQ_PINLOC_8),
      .PORT_MEM_DQ_PINLOC_9 (PORT_MEM_DQ_PINLOC_9),
      .PORT_MEM_DQ_PINLOC_10 (PORT_MEM_DQ_PINLOC_10),
      .PORT_MEM_DQ_PINLOC_11 (PORT_MEM_DQ_PINLOC_11),
      .PORT_MEM_DQ_PINLOC_12 (PORT_MEM_DQ_PINLOC_12),
      .PORT_MEM_DQ_PINLOC_13 (PORT_MEM_DQ_PINLOC_13),
      .PORT_MEM_DQ_PINLOC_14 (PORT_MEM_DQ_PINLOC_14),
      .PORT_MEM_DQ_PINLOC_15 (PORT_MEM_DQ_PINLOC_15),
      .PORT_MEM_DQ_PINLOC_16 (PORT_MEM_DQ_PINLOC_16),
      .PORT_MEM_DQ_PINLOC_17 (PORT_MEM_DQ_PINLOC_17),
      .PORT_MEM_DQ_PINLOC_18 (PORT_MEM_DQ_PINLOC_18),
      .PORT_MEM_DQ_PINLOC_19 (PORT_MEM_DQ_PINLOC_19),
      .PORT_MEM_DQ_PINLOC_20 (PORT_MEM_DQ_PINLOC_20),
      .PORT_MEM_DQ_PINLOC_21 (PORT_MEM_DQ_PINLOC_21),
      .PORT_MEM_DQ_PINLOC_22 (PORT_MEM_DQ_PINLOC_22),
      .PORT_MEM_DQ_PINLOC_23 (PORT_MEM_DQ_PINLOC_23),
      .PORT_MEM_DQ_PINLOC_24 (PORT_MEM_DQ_PINLOC_24),
      .PORT_MEM_DQ_PINLOC_25 (PORT_MEM_DQ_PINLOC_25),
      .PORT_MEM_DQ_PINLOC_26 (PORT_MEM_DQ_PINLOC_26),
      .PORT_MEM_DQ_PINLOC_27 (PORT_MEM_DQ_PINLOC_27),
      .PORT_MEM_DQ_PINLOC_28 (PORT_MEM_DQ_PINLOC_28),
      .PORT_MEM_DQ_PINLOC_29 (PORT_MEM_DQ_PINLOC_29),
      .PORT_MEM_DQ_PINLOC_30 (PORT_MEM_DQ_PINLOC_30),
      .PORT_MEM_DQ_PINLOC_31 (PORT_MEM_DQ_PINLOC_31),
      .PORT_MEM_DQ_PINLOC_32 (PORT_MEM_DQ_PINLOC_32),
      .PORT_MEM_DQ_PINLOC_33 (PORT_MEM_DQ_PINLOC_33),
      .PORT_MEM_DQ_PINLOC_34 (PORT_MEM_DQ_PINLOC_34),
      .PORT_MEM_DQ_PINLOC_35 (PORT_MEM_DQ_PINLOC_35),
      .PORT_MEM_DQ_PINLOC_36 (PORT_MEM_DQ_PINLOC_36),
      .PORT_MEM_DQ_PINLOC_37 (PORT_MEM_DQ_PINLOC_37),
      .PORT_MEM_DQ_PINLOC_38 (PORT_MEM_DQ_PINLOC_38),
      .PORT_MEM_DQ_PINLOC_39 (PORT_MEM_DQ_PINLOC_39),
      .PORT_MEM_DQ_PINLOC_40 (PORT_MEM_DQ_PINLOC_40),
      .PORT_MEM_DQ_PINLOC_41 (PORT_MEM_DQ_PINLOC_41),
      .PORT_MEM_DQ_PINLOC_42 (PORT_MEM_DQ_PINLOC_42),
      .PORT_MEM_DQ_PINLOC_43 (PORT_MEM_DQ_PINLOC_43),
      .PORT_MEM_DQ_PINLOC_44 (PORT_MEM_DQ_PINLOC_44),
      .PORT_MEM_DQ_PINLOC_45 (PORT_MEM_DQ_PINLOC_45),
      .PORT_MEM_DQ_PINLOC_46 (PORT_MEM_DQ_PINLOC_46),
      .PORT_MEM_DQ_PINLOC_47 (PORT_MEM_DQ_PINLOC_47),
      .PORT_MEM_DQ_PINLOC_48 (PORT_MEM_DQ_PINLOC_48),
      .PORT_MEM_DQ_PINLOC_AUTOGEN_WCNT (PORT_MEM_DQ_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DBI_N_WIDTH (PORT_MEM_DBI_N_WIDTH),
      .PORT_MEM_DBI_N_PINLOC_0 (PORT_MEM_DBI_N_PINLOC_0),
      .PORT_MEM_DBI_N_PINLOC_1 (PORT_MEM_DBI_N_PINLOC_1),
      .PORT_MEM_DBI_N_PINLOC_2 (PORT_MEM_DBI_N_PINLOC_2),
      .PORT_MEM_DBI_N_PINLOC_3 (PORT_MEM_DBI_N_PINLOC_3),
      .PORT_MEM_DBI_N_PINLOC_4 (PORT_MEM_DBI_N_PINLOC_4),
      .PORT_MEM_DBI_N_PINLOC_5 (PORT_MEM_DBI_N_PINLOC_5),
      .PORT_MEM_DBI_N_PINLOC_6 (PORT_MEM_DBI_N_PINLOC_6),
      .PORT_MEM_DBI_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_DBI_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DQA_WIDTH (PORT_MEM_DQA_WIDTH),
      .PORT_MEM_DQA_PINLOC_0 (PORT_MEM_DQA_PINLOC_0),
      .PORT_MEM_DQA_PINLOC_1 (PORT_MEM_DQA_PINLOC_1),
      .PORT_MEM_DQA_PINLOC_2 (PORT_MEM_DQA_PINLOC_2),
      .PORT_MEM_DQA_PINLOC_3 (PORT_MEM_DQA_PINLOC_3),
      .PORT_MEM_DQA_PINLOC_4 (PORT_MEM_DQA_PINLOC_4),
      .PORT_MEM_DQA_PINLOC_5 (PORT_MEM_DQA_PINLOC_5),
      .PORT_MEM_DQA_PINLOC_6 (PORT_MEM_DQA_PINLOC_6),
      .PORT_MEM_DQA_PINLOC_7 (PORT_MEM_DQA_PINLOC_7),
      .PORT_MEM_DQA_PINLOC_8 (PORT_MEM_DQA_PINLOC_8),
      .PORT_MEM_DQA_PINLOC_9 (PORT_MEM_DQA_PINLOC_9),
      .PORT_MEM_DQA_PINLOC_10 (PORT_MEM_DQA_PINLOC_10),
      .PORT_MEM_DQA_PINLOC_11 (PORT_MEM_DQA_PINLOC_11),
      .PORT_MEM_DQA_PINLOC_12 (PORT_MEM_DQA_PINLOC_12),
      .PORT_MEM_DQA_PINLOC_13 (PORT_MEM_DQA_PINLOC_13),
      .PORT_MEM_DQA_PINLOC_14 (PORT_MEM_DQA_PINLOC_14),
      .PORT_MEM_DQA_PINLOC_15 (PORT_MEM_DQA_PINLOC_15),
      .PORT_MEM_DQA_PINLOC_16 (PORT_MEM_DQA_PINLOC_16),
      .PORT_MEM_DQA_PINLOC_17 (PORT_MEM_DQA_PINLOC_17),
      .PORT_MEM_DQA_PINLOC_18 (PORT_MEM_DQA_PINLOC_18),
      .PORT_MEM_DQA_PINLOC_19 (PORT_MEM_DQA_PINLOC_19),
      .PORT_MEM_DQA_PINLOC_20 (PORT_MEM_DQA_PINLOC_20),
      .PORT_MEM_DQA_PINLOC_21 (PORT_MEM_DQA_PINLOC_21),
      .PORT_MEM_DQA_PINLOC_22 (PORT_MEM_DQA_PINLOC_22),
      .PORT_MEM_DQA_PINLOC_23 (PORT_MEM_DQA_PINLOC_23),
      .PORT_MEM_DQA_PINLOC_24 (PORT_MEM_DQA_PINLOC_24),
      .PORT_MEM_DQA_PINLOC_25 (PORT_MEM_DQA_PINLOC_25),
      .PORT_MEM_DQA_PINLOC_26 (PORT_MEM_DQA_PINLOC_26),
      .PORT_MEM_DQA_PINLOC_27 (PORT_MEM_DQA_PINLOC_27),
      .PORT_MEM_DQA_PINLOC_28 (PORT_MEM_DQA_PINLOC_28),
      .PORT_MEM_DQA_PINLOC_29 (PORT_MEM_DQA_PINLOC_29),
      .PORT_MEM_DQA_PINLOC_30 (PORT_MEM_DQA_PINLOC_30),
      .PORT_MEM_DQA_PINLOC_31 (PORT_MEM_DQA_PINLOC_31),
      .PORT_MEM_DQA_PINLOC_32 (PORT_MEM_DQA_PINLOC_32),
      .PORT_MEM_DQA_PINLOC_33 (PORT_MEM_DQA_PINLOC_33),
      .PORT_MEM_DQA_PINLOC_34 (PORT_MEM_DQA_PINLOC_34),
      .PORT_MEM_DQA_PINLOC_35 (PORT_MEM_DQA_PINLOC_35),
      .PORT_MEM_DQA_PINLOC_36 (PORT_MEM_DQA_PINLOC_36),
      .PORT_MEM_DQA_PINLOC_37 (PORT_MEM_DQA_PINLOC_37),
      .PORT_MEM_DQA_PINLOC_38 (PORT_MEM_DQA_PINLOC_38),
      .PORT_MEM_DQA_PINLOC_39 (PORT_MEM_DQA_PINLOC_39),
      .PORT_MEM_DQA_PINLOC_40 (PORT_MEM_DQA_PINLOC_40),
      .PORT_MEM_DQA_PINLOC_41 (PORT_MEM_DQA_PINLOC_41),
      .PORT_MEM_DQA_PINLOC_42 (PORT_MEM_DQA_PINLOC_42),
      .PORT_MEM_DQA_PINLOC_43 (PORT_MEM_DQA_PINLOC_43),
      .PORT_MEM_DQA_PINLOC_44 (PORT_MEM_DQA_PINLOC_44),
      .PORT_MEM_DQA_PINLOC_45 (PORT_MEM_DQA_PINLOC_45),
      .PORT_MEM_DQA_PINLOC_46 (PORT_MEM_DQA_PINLOC_46),
      .PORT_MEM_DQA_PINLOC_47 (PORT_MEM_DQA_PINLOC_47),
      .PORT_MEM_DQA_PINLOC_48 (PORT_MEM_DQA_PINLOC_48),
      .PORT_MEM_DQA_PINLOC_AUTOGEN_WCNT (PORT_MEM_DQA_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DQB_WIDTH (PORT_MEM_DQB_WIDTH),
      .PORT_MEM_DQB_PINLOC_0 (PORT_MEM_DQB_PINLOC_0),
      .PORT_MEM_DQB_PINLOC_1 (PORT_MEM_DQB_PINLOC_1),
      .PORT_MEM_DQB_PINLOC_2 (PORT_MEM_DQB_PINLOC_2),
      .PORT_MEM_DQB_PINLOC_3 (PORT_MEM_DQB_PINLOC_3),
      .PORT_MEM_DQB_PINLOC_4 (PORT_MEM_DQB_PINLOC_4),
      .PORT_MEM_DQB_PINLOC_5 (PORT_MEM_DQB_PINLOC_5),
      .PORT_MEM_DQB_PINLOC_6 (PORT_MEM_DQB_PINLOC_6),
      .PORT_MEM_DQB_PINLOC_7 (PORT_MEM_DQB_PINLOC_7),
      .PORT_MEM_DQB_PINLOC_8 (PORT_MEM_DQB_PINLOC_8),
      .PORT_MEM_DQB_PINLOC_9 (PORT_MEM_DQB_PINLOC_9),
      .PORT_MEM_DQB_PINLOC_10 (PORT_MEM_DQB_PINLOC_10),
      .PORT_MEM_DQB_PINLOC_11 (PORT_MEM_DQB_PINLOC_11),
      .PORT_MEM_DQB_PINLOC_12 (PORT_MEM_DQB_PINLOC_12),
      .PORT_MEM_DQB_PINLOC_13 (PORT_MEM_DQB_PINLOC_13),
      .PORT_MEM_DQB_PINLOC_14 (PORT_MEM_DQB_PINLOC_14),
      .PORT_MEM_DQB_PINLOC_15 (PORT_MEM_DQB_PINLOC_15),
      .PORT_MEM_DQB_PINLOC_16 (PORT_MEM_DQB_PINLOC_16),
      .PORT_MEM_DQB_PINLOC_17 (PORT_MEM_DQB_PINLOC_17),
      .PORT_MEM_DQB_PINLOC_18 (PORT_MEM_DQB_PINLOC_18),
      .PORT_MEM_DQB_PINLOC_19 (PORT_MEM_DQB_PINLOC_19),
      .PORT_MEM_DQB_PINLOC_20 (PORT_MEM_DQB_PINLOC_20),
      .PORT_MEM_DQB_PINLOC_21 (PORT_MEM_DQB_PINLOC_21),
      .PORT_MEM_DQB_PINLOC_22 (PORT_MEM_DQB_PINLOC_22),
      .PORT_MEM_DQB_PINLOC_23 (PORT_MEM_DQB_PINLOC_23),
      .PORT_MEM_DQB_PINLOC_24 (PORT_MEM_DQB_PINLOC_24),
      .PORT_MEM_DQB_PINLOC_25 (PORT_MEM_DQB_PINLOC_25),
      .PORT_MEM_DQB_PINLOC_26 (PORT_MEM_DQB_PINLOC_26),
      .PORT_MEM_DQB_PINLOC_27 (PORT_MEM_DQB_PINLOC_27),
      .PORT_MEM_DQB_PINLOC_28 (PORT_MEM_DQB_PINLOC_28),
      .PORT_MEM_DQB_PINLOC_29 (PORT_MEM_DQB_PINLOC_29),
      .PORT_MEM_DQB_PINLOC_30 (PORT_MEM_DQB_PINLOC_30),
      .PORT_MEM_DQB_PINLOC_31 (PORT_MEM_DQB_PINLOC_31),
      .PORT_MEM_DQB_PINLOC_32 (PORT_MEM_DQB_PINLOC_32),
      .PORT_MEM_DQB_PINLOC_33 (PORT_MEM_DQB_PINLOC_33),
      .PORT_MEM_DQB_PINLOC_34 (PORT_MEM_DQB_PINLOC_34),
      .PORT_MEM_DQB_PINLOC_35 (PORT_MEM_DQB_PINLOC_35),
      .PORT_MEM_DQB_PINLOC_36 (PORT_MEM_DQB_PINLOC_36),
      .PORT_MEM_DQB_PINLOC_37 (PORT_MEM_DQB_PINLOC_37),
      .PORT_MEM_DQB_PINLOC_38 (PORT_MEM_DQB_PINLOC_38),
      .PORT_MEM_DQB_PINLOC_39 (PORT_MEM_DQB_PINLOC_39),
      .PORT_MEM_DQB_PINLOC_40 (PORT_MEM_DQB_PINLOC_40),
      .PORT_MEM_DQB_PINLOC_41 (PORT_MEM_DQB_PINLOC_41),
      .PORT_MEM_DQB_PINLOC_42 (PORT_MEM_DQB_PINLOC_42),
      .PORT_MEM_DQB_PINLOC_43 (PORT_MEM_DQB_PINLOC_43),
      .PORT_MEM_DQB_PINLOC_44 (PORT_MEM_DQB_PINLOC_44),
      .PORT_MEM_DQB_PINLOC_45 (PORT_MEM_DQB_PINLOC_45),
      .PORT_MEM_DQB_PINLOC_46 (PORT_MEM_DQB_PINLOC_46),
      .PORT_MEM_DQB_PINLOC_47 (PORT_MEM_DQB_PINLOC_47),
      .PORT_MEM_DQB_PINLOC_48 (PORT_MEM_DQB_PINLOC_48),
      .PORT_MEM_DQB_PINLOC_AUTOGEN_WCNT (PORT_MEM_DQB_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DINVA_WIDTH (PORT_MEM_DINVA_WIDTH),
      .PORT_MEM_DINVA_PINLOC_0 (PORT_MEM_DINVA_PINLOC_0),
      .PORT_MEM_DINVA_PINLOC_1 (PORT_MEM_DINVA_PINLOC_1),
      .PORT_MEM_DINVA_PINLOC_2 (PORT_MEM_DINVA_PINLOC_2),
      .PORT_MEM_DINVA_PINLOC_AUTOGEN_WCNT (PORT_MEM_DINVA_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DINVB_WIDTH (PORT_MEM_DINVB_WIDTH),
      .PORT_MEM_DINVB_PINLOC_0 (PORT_MEM_DINVB_PINLOC_0),
      .PORT_MEM_DINVB_PINLOC_1 (PORT_MEM_DINVB_PINLOC_1),
      .PORT_MEM_DINVB_PINLOC_2 (PORT_MEM_DINVB_PINLOC_2),
      .PORT_MEM_DINVB_PINLOC_AUTOGEN_WCNT (PORT_MEM_DINVB_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_Q_WIDTH (PORT_MEM_Q_WIDTH),
      .PORT_MEM_Q_PINLOC_0 (PORT_MEM_Q_PINLOC_0),
      .PORT_MEM_Q_PINLOC_1 (PORT_MEM_Q_PINLOC_1),
      .PORT_MEM_Q_PINLOC_2 (PORT_MEM_Q_PINLOC_2),
      .PORT_MEM_Q_PINLOC_3 (PORT_MEM_Q_PINLOC_3),
      .PORT_MEM_Q_PINLOC_4 (PORT_MEM_Q_PINLOC_4),
      .PORT_MEM_Q_PINLOC_5 (PORT_MEM_Q_PINLOC_5),
      .PORT_MEM_Q_PINLOC_6 (PORT_MEM_Q_PINLOC_6),
      .PORT_MEM_Q_PINLOC_7 (PORT_MEM_Q_PINLOC_7),
      .PORT_MEM_Q_PINLOC_8 (PORT_MEM_Q_PINLOC_8),
      .PORT_MEM_Q_PINLOC_9 (PORT_MEM_Q_PINLOC_9),
      .PORT_MEM_Q_PINLOC_10 (PORT_MEM_Q_PINLOC_10),
      .PORT_MEM_Q_PINLOC_11 (PORT_MEM_Q_PINLOC_11),
      .PORT_MEM_Q_PINLOC_12 (PORT_MEM_Q_PINLOC_12),
      .PORT_MEM_Q_PINLOC_13 (PORT_MEM_Q_PINLOC_13),
      .PORT_MEM_Q_PINLOC_14 (PORT_MEM_Q_PINLOC_14),
      .PORT_MEM_Q_PINLOC_15 (PORT_MEM_Q_PINLOC_15),
      .PORT_MEM_Q_PINLOC_16 (PORT_MEM_Q_PINLOC_16),
      .PORT_MEM_Q_PINLOC_17 (PORT_MEM_Q_PINLOC_17),
      .PORT_MEM_Q_PINLOC_18 (PORT_MEM_Q_PINLOC_18),
      .PORT_MEM_Q_PINLOC_19 (PORT_MEM_Q_PINLOC_19),
      .PORT_MEM_Q_PINLOC_20 (PORT_MEM_Q_PINLOC_20),
      .PORT_MEM_Q_PINLOC_21 (PORT_MEM_Q_PINLOC_21),
      .PORT_MEM_Q_PINLOC_22 (PORT_MEM_Q_PINLOC_22),
      .PORT_MEM_Q_PINLOC_23 (PORT_MEM_Q_PINLOC_23),
      .PORT_MEM_Q_PINLOC_24 (PORT_MEM_Q_PINLOC_24),
      .PORT_MEM_Q_PINLOC_25 (PORT_MEM_Q_PINLOC_25),
      .PORT_MEM_Q_PINLOC_26 (PORT_MEM_Q_PINLOC_26),
      .PORT_MEM_Q_PINLOC_27 (PORT_MEM_Q_PINLOC_27),
      .PORT_MEM_Q_PINLOC_28 (PORT_MEM_Q_PINLOC_28),
      .PORT_MEM_Q_PINLOC_29 (PORT_MEM_Q_PINLOC_29),
      .PORT_MEM_Q_PINLOC_30 (PORT_MEM_Q_PINLOC_30),
      .PORT_MEM_Q_PINLOC_31 (PORT_MEM_Q_PINLOC_31),
      .PORT_MEM_Q_PINLOC_32 (PORT_MEM_Q_PINLOC_32),
      .PORT_MEM_Q_PINLOC_33 (PORT_MEM_Q_PINLOC_33),
      .PORT_MEM_Q_PINLOC_34 (PORT_MEM_Q_PINLOC_34),
      .PORT_MEM_Q_PINLOC_35 (PORT_MEM_Q_PINLOC_35),
      .PORT_MEM_Q_PINLOC_36 (PORT_MEM_Q_PINLOC_36),
      .PORT_MEM_Q_PINLOC_37 (PORT_MEM_Q_PINLOC_37),
      .PORT_MEM_Q_PINLOC_38 (PORT_MEM_Q_PINLOC_38),
      .PORT_MEM_Q_PINLOC_39 (PORT_MEM_Q_PINLOC_39),
      .PORT_MEM_Q_PINLOC_40 (PORT_MEM_Q_PINLOC_40),
      .PORT_MEM_Q_PINLOC_41 (PORT_MEM_Q_PINLOC_41),
      .PORT_MEM_Q_PINLOC_42 (PORT_MEM_Q_PINLOC_42),
      .PORT_MEM_Q_PINLOC_43 (PORT_MEM_Q_PINLOC_43),
      .PORT_MEM_Q_PINLOC_44 (PORT_MEM_Q_PINLOC_44),
      .PORT_MEM_Q_PINLOC_45 (PORT_MEM_Q_PINLOC_45),
      .PORT_MEM_Q_PINLOC_46 (PORT_MEM_Q_PINLOC_46),
      .PORT_MEM_Q_PINLOC_47 (PORT_MEM_Q_PINLOC_47),
      .PORT_MEM_Q_PINLOC_48 (PORT_MEM_Q_PINLOC_48),
      .PORT_MEM_Q_PINLOC_AUTOGEN_WCNT (PORT_MEM_Q_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DQS_WIDTH (PORT_MEM_DQS_WIDTH),
      .PORT_MEM_DQS_PINLOC_0 (PORT_MEM_DQS_PINLOC_0),
      .PORT_MEM_DQS_PINLOC_1 (PORT_MEM_DQS_PINLOC_1),
      .PORT_MEM_DQS_PINLOC_2 (PORT_MEM_DQS_PINLOC_2),
      .PORT_MEM_DQS_PINLOC_3 (PORT_MEM_DQS_PINLOC_3),
      .PORT_MEM_DQS_PINLOC_4 (PORT_MEM_DQS_PINLOC_4),
      .PORT_MEM_DQS_PINLOC_5 (PORT_MEM_DQS_PINLOC_5),
      .PORT_MEM_DQS_PINLOC_6 (PORT_MEM_DQS_PINLOC_6),
      .PORT_MEM_DQS_PINLOC_7 (PORT_MEM_DQS_PINLOC_7),
      .PORT_MEM_DQS_PINLOC_8 (PORT_MEM_DQS_PINLOC_8),
      .PORT_MEM_DQS_PINLOC_9 (PORT_MEM_DQS_PINLOC_9),
      .PORT_MEM_DQS_PINLOC_10 (PORT_MEM_DQS_PINLOC_10),
      .PORT_MEM_DQS_PINLOC_11 (PORT_MEM_DQS_PINLOC_11),
      .PORT_MEM_DQS_PINLOC_12 (PORT_MEM_DQS_PINLOC_12),
      .PORT_MEM_DQS_PINLOC_AUTOGEN_WCNT (PORT_MEM_DQS_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_DQS_N_WIDTH (PORT_MEM_DQS_N_WIDTH),
      .PORT_MEM_DQS_N_PINLOC_0 (PORT_MEM_DQS_N_PINLOC_0),
      .PORT_MEM_DQS_N_PINLOC_1 (PORT_MEM_DQS_N_PINLOC_1),
      .PORT_MEM_DQS_N_PINLOC_2 (PORT_MEM_DQS_N_PINLOC_2),
      .PORT_MEM_DQS_N_PINLOC_3 (PORT_MEM_DQS_N_PINLOC_3),
      .PORT_MEM_DQS_N_PINLOC_4 (PORT_MEM_DQS_N_PINLOC_4),
      .PORT_MEM_DQS_N_PINLOC_5 (PORT_MEM_DQS_N_PINLOC_5),
      .PORT_MEM_DQS_N_PINLOC_6 (PORT_MEM_DQS_N_PINLOC_6),
      .PORT_MEM_DQS_N_PINLOC_7 (PORT_MEM_DQS_N_PINLOC_7),
      .PORT_MEM_DQS_N_PINLOC_8 (PORT_MEM_DQS_N_PINLOC_8),
      .PORT_MEM_DQS_N_PINLOC_9 (PORT_MEM_DQS_N_PINLOC_9),
      .PORT_MEM_DQS_N_PINLOC_10 (PORT_MEM_DQS_N_PINLOC_10),
      .PORT_MEM_DQS_N_PINLOC_11 (PORT_MEM_DQS_N_PINLOC_11),
      .PORT_MEM_DQS_N_PINLOC_12 (PORT_MEM_DQS_N_PINLOC_12),
      .PORT_MEM_DQS_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_DQS_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_QK_WIDTH (PORT_MEM_QK_WIDTH),
      .PORT_MEM_QK_PINLOC_0 (PORT_MEM_QK_PINLOC_0),
      .PORT_MEM_QK_PINLOC_1 (PORT_MEM_QK_PINLOC_1),
      .PORT_MEM_QK_PINLOC_2 (PORT_MEM_QK_PINLOC_2),
      .PORT_MEM_QK_PINLOC_3 (PORT_MEM_QK_PINLOC_3),
      .PORT_MEM_QK_PINLOC_4 (PORT_MEM_QK_PINLOC_4),
      .PORT_MEM_QK_PINLOC_5 (PORT_MEM_QK_PINLOC_5),
      .PORT_MEM_QK_PINLOC_AUTOGEN_WCNT (PORT_MEM_QK_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_QK_N_WIDTH (PORT_MEM_QK_N_WIDTH),
      .PORT_MEM_QK_N_PINLOC_0 (PORT_MEM_QK_N_PINLOC_0),
      .PORT_MEM_QK_N_PINLOC_1 (PORT_MEM_QK_N_PINLOC_1),
      .PORT_MEM_QK_N_PINLOC_2 (PORT_MEM_QK_N_PINLOC_2),
      .PORT_MEM_QK_N_PINLOC_3 (PORT_MEM_QK_N_PINLOC_3),
      .PORT_MEM_QK_N_PINLOC_4 (PORT_MEM_QK_N_PINLOC_4),
      .PORT_MEM_QK_N_PINLOC_5 (PORT_MEM_QK_N_PINLOC_5),
      .PORT_MEM_QK_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_QK_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_QKA_WIDTH (PORT_MEM_QKA_WIDTH),
      .PORT_MEM_QKA_PINLOC_0 (PORT_MEM_QKA_PINLOC_0),
      .PORT_MEM_QKA_PINLOC_1 (PORT_MEM_QKA_PINLOC_1),
      .PORT_MEM_QKA_PINLOC_2 (PORT_MEM_QKA_PINLOC_2),
      .PORT_MEM_QKA_PINLOC_3 (PORT_MEM_QKA_PINLOC_3),
      .PORT_MEM_QKA_PINLOC_4 (PORT_MEM_QKA_PINLOC_4),
      .PORT_MEM_QKA_PINLOC_5 (PORT_MEM_QKA_PINLOC_5),
      .PORT_MEM_QKA_PINLOC_AUTOGEN_WCNT (PORT_MEM_QKA_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_QKA_N_WIDTH (PORT_MEM_QKA_N_WIDTH),
      .PORT_MEM_QKA_N_PINLOC_0 (PORT_MEM_QKA_N_PINLOC_0),
      .PORT_MEM_QKA_N_PINLOC_1 (PORT_MEM_QKA_N_PINLOC_1),
      .PORT_MEM_QKA_N_PINLOC_2 (PORT_MEM_QKA_N_PINLOC_2),
      .PORT_MEM_QKA_N_PINLOC_3 (PORT_MEM_QKA_N_PINLOC_3),
      .PORT_MEM_QKA_N_PINLOC_4 (PORT_MEM_QKA_N_PINLOC_4),
      .PORT_MEM_QKA_N_PINLOC_5 (PORT_MEM_QKA_N_PINLOC_5),
      .PORT_MEM_QKA_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_QKA_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_QKB_WIDTH (PORT_MEM_QKB_WIDTH),
      .PORT_MEM_QKB_PINLOC_0 (PORT_MEM_QKB_PINLOC_0),
      .PORT_MEM_QKB_PINLOC_1 (PORT_MEM_QKB_PINLOC_1),
      .PORT_MEM_QKB_PINLOC_2 (PORT_MEM_QKB_PINLOC_2),
      .PORT_MEM_QKB_PINLOC_3 (PORT_MEM_QKB_PINLOC_3),
      .PORT_MEM_QKB_PINLOC_4 (PORT_MEM_QKB_PINLOC_4),
      .PORT_MEM_QKB_PINLOC_5 (PORT_MEM_QKB_PINLOC_5),
      .PORT_MEM_QKB_PINLOC_AUTOGEN_WCNT (PORT_MEM_QKB_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_QKB_N_WIDTH (PORT_MEM_QKB_N_WIDTH),
      .PORT_MEM_QKB_N_PINLOC_0 (PORT_MEM_QKB_N_PINLOC_0),
      .PORT_MEM_QKB_N_PINLOC_1 (PORT_MEM_QKB_N_PINLOC_1),
      .PORT_MEM_QKB_N_PINLOC_2 (PORT_MEM_QKB_N_PINLOC_2),
      .PORT_MEM_QKB_N_PINLOC_3 (PORT_MEM_QKB_N_PINLOC_3),
      .PORT_MEM_QKB_N_PINLOC_4 (PORT_MEM_QKB_N_PINLOC_4),
      .PORT_MEM_QKB_N_PINLOC_5 (PORT_MEM_QKB_N_PINLOC_5),
      .PORT_MEM_QKB_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_QKB_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CQ_WIDTH (PORT_MEM_CQ_WIDTH),
      .PORT_MEM_CQ_PINLOC_0 (PORT_MEM_CQ_PINLOC_0),
      .PORT_MEM_CQ_PINLOC_1 (PORT_MEM_CQ_PINLOC_1),
      .PORT_MEM_CQ_PINLOC_AUTOGEN_WCNT (PORT_MEM_CQ_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_CQ_N_WIDTH (PORT_MEM_CQ_N_WIDTH),
      .PORT_MEM_CQ_N_PINLOC_0 (PORT_MEM_CQ_N_PINLOC_0),
      .PORT_MEM_CQ_N_PINLOC_1 (PORT_MEM_CQ_N_PINLOC_1),
      .PORT_MEM_CQ_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_CQ_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_ALERT_N_WIDTH (PORT_MEM_ALERT_N_WIDTH),
      .PORT_MEM_ALERT_N_PINLOC_0 (PORT_MEM_ALERT_N_PINLOC_0),
      .PORT_MEM_ALERT_N_PINLOC_1 (PORT_MEM_ALERT_N_PINLOC_1),
      .PORT_MEM_ALERT_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_ALERT_N_PINLOC_AUTOGEN_WCNT),
      .PORT_MEM_PE_N_WIDTH (PORT_MEM_PE_N_WIDTH),
      .PORT_MEM_PE_N_PINLOC_0 (PORT_MEM_PE_N_PINLOC_0),
      .PORT_MEM_PE_N_PINLOC_1 (PORT_MEM_PE_N_PINLOC_1),
      .PORT_MEM_PE_N_PINLOC_AUTOGEN_WCNT (PORT_MEM_PE_N_PINLOC_AUTOGEN_WCNT),
      .PORT_CLKS_SHARING_MASTER_OUT_WIDTH (PORT_CLKS_SHARING_MASTER_OUT_WIDTH),
      .PORT_CLKS_SHARING_SLAVE_IN_WIDTH (PORT_CLKS_SHARING_SLAVE_IN_WIDTH),
      .PORT_AFI_RLAT_WIDTH (PORT_AFI_RLAT_WIDTH),
      .PORT_AFI_WLAT_WIDTH (PORT_AFI_WLAT_WIDTH),
      .PORT_AFI_SEQ_BUSY_WIDTH (PORT_AFI_SEQ_BUSY_WIDTH),
      .PORT_AFI_ADDR_WIDTH (PORT_AFI_ADDR_WIDTH),
      .PORT_AFI_BA_WIDTH (PORT_AFI_BA_WIDTH),
      .PORT_AFI_BG_WIDTH (PORT_AFI_BG_WIDTH),
      .PORT_AFI_C_WIDTH (PORT_AFI_C_WIDTH),
      .PORT_AFI_CKE_WIDTH (PORT_AFI_CKE_WIDTH),
      .PORT_AFI_CS_N_WIDTH (PORT_AFI_CS_N_WIDTH),
      .PORT_AFI_RM_WIDTH (PORT_AFI_RM_WIDTH),
      .PORT_AFI_ODT_WIDTH (PORT_AFI_ODT_WIDTH),
      .PORT_AFI_RAS_N_WIDTH (PORT_AFI_RAS_N_WIDTH),
      .PORT_AFI_CAS_N_WIDTH (PORT_AFI_CAS_N_WIDTH),
      .PORT_AFI_WE_N_WIDTH (PORT_AFI_WE_N_WIDTH),
      .PORT_AFI_RST_N_WIDTH (PORT_AFI_RST_N_WIDTH),
      .PORT_AFI_ACT_N_WIDTH (PORT_AFI_ACT_N_WIDTH),
      .PORT_AFI_PAR_WIDTH (PORT_AFI_PAR_WIDTH),
      .PORT_AFI_CA_WIDTH (PORT_AFI_CA_WIDTH),
      .PORT_AFI_REF_N_WIDTH (PORT_AFI_REF_N_WIDTH),
      .PORT_AFI_WPS_N_WIDTH (PORT_AFI_WPS_N_WIDTH),
      .PORT_AFI_RPS_N_WIDTH (PORT_AFI_RPS_N_WIDTH),
      .PORT_AFI_DOFF_N_WIDTH (PORT_AFI_DOFF_N_WIDTH),
      .PORT_AFI_LD_N_WIDTH (PORT_AFI_LD_N_WIDTH),
      .PORT_AFI_RW_N_WIDTH (PORT_AFI_RW_N_WIDTH),
      .PORT_AFI_LBK0_N_WIDTH (PORT_AFI_LBK0_N_WIDTH),
      .PORT_AFI_LBK1_N_WIDTH (PORT_AFI_LBK1_N_WIDTH),
      .PORT_AFI_CFG_N_WIDTH (PORT_AFI_CFG_N_WIDTH),
      .PORT_AFI_AP_WIDTH (PORT_AFI_AP_WIDTH),
      .PORT_AFI_AINV_WIDTH (PORT_AFI_AINV_WIDTH),
      .PORT_AFI_DM_WIDTH (PORT_AFI_DM_WIDTH),
      .PORT_AFI_DM_N_WIDTH (PORT_AFI_DM_N_WIDTH),
      .PORT_AFI_BWS_N_WIDTH (PORT_AFI_BWS_N_WIDTH),
      .PORT_AFI_RDATA_DBI_N_WIDTH (PORT_AFI_RDATA_DBI_N_WIDTH),
      .PORT_AFI_WDATA_DBI_N_WIDTH (PORT_AFI_WDATA_DBI_N_WIDTH),
      .PORT_AFI_RDATA_DINV_WIDTH (PORT_AFI_RDATA_DINV_WIDTH),
      .PORT_AFI_WDATA_DINV_WIDTH (PORT_AFI_WDATA_DINV_WIDTH),
      .PORT_AFI_DQS_BURST_WIDTH (PORT_AFI_DQS_BURST_WIDTH),
      .PORT_AFI_WDATA_VALID_WIDTH (PORT_AFI_WDATA_VALID_WIDTH),
      .PORT_AFI_WDATA_WIDTH (PORT_AFI_WDATA_WIDTH),
      .PORT_AFI_RDATA_EN_FULL_WIDTH (PORT_AFI_RDATA_EN_FULL_WIDTH),
      .PORT_AFI_RDATA_WIDTH (PORT_AFI_RDATA_WIDTH),
      .PORT_AFI_RDATA_VALID_WIDTH (PORT_AFI_RDATA_VALID_WIDTH),
      .PORT_AFI_RRANK_WIDTH (PORT_AFI_RRANK_WIDTH),
      .PORT_AFI_WRANK_WIDTH (PORT_AFI_WRANK_WIDTH),
      .PORT_AFI_ALERT_N_WIDTH (PORT_AFI_ALERT_N_WIDTH),
      .PORT_AFI_PE_N_WIDTH (PORT_AFI_PE_N_WIDTH),
      .PORT_CTRL_AST_CMD_DATA_WIDTH (PORT_CTRL_AST_CMD_DATA_WIDTH),
      .PORT_CTRL_AST_WR_DATA_WIDTH (PORT_CTRL_AST_WR_DATA_WIDTH),
      .PORT_CTRL_AST_RD_DATA_WIDTH (PORT_CTRL_AST_RD_DATA_WIDTH),
      .PORT_CTRL_AMM_ADDRESS_WIDTH (PORT_CTRL_AMM_ADDRESS_WIDTH),
      .PORT_CTRL_AMM_RDATA_WIDTH (PORT_CTRL_AMM_RDATA_WIDTH),
      .PORT_CTRL_AMM_WDATA_WIDTH (PORT_CTRL_AMM_WDATA_WIDTH),
      .PORT_CTRL_AMM_BCOUNT_WIDTH (PORT_CTRL_AMM_BCOUNT_WIDTH),
      .PORT_CTRL_AMM_BYTEEN_WIDTH (PORT_CTRL_AMM_BYTEEN_WIDTH),
      .PORT_CTRL_USER_REFRESH_REQ_WIDTH (PORT_CTRL_USER_REFRESH_REQ_WIDTH),
      .PORT_CTRL_USER_REFRESH_BANK_WIDTH (PORT_CTRL_USER_REFRESH_BANK_WIDTH),
      .PORT_CTRL_SELF_REFRESH_REQ_WIDTH (PORT_CTRL_SELF_REFRESH_REQ_WIDTH),
      .PORT_CTRL_ECC_WRITE_INFO_WIDTH (PORT_CTRL_ECC_WRITE_INFO_WIDTH),
      .PORT_CTRL_ECC_RDATA_ID_WIDTH (PORT_CTRL_ECC_RDATA_ID_WIDTH),
      .PORT_CTRL_ECC_READ_INFO_WIDTH (PORT_CTRL_ECC_READ_INFO_WIDTH),
      .PORT_CTRL_ECC_CMD_INFO_WIDTH (PORT_CTRL_ECC_CMD_INFO_WIDTH),
      .PORT_CTRL_ECC_WB_POINTER_WIDTH (PORT_CTRL_ECC_WB_POINTER_WIDTH),
      .PORT_CTRL_MMR_SLAVE_ADDRESS_WIDTH (PORT_CTRL_MMR_SLAVE_ADDRESS_WIDTH),
      .PORT_CTRL_MMR_SLAVE_RDATA_WIDTH (PORT_CTRL_MMR_SLAVE_RDATA_WIDTH),
      .PORT_CTRL_MMR_SLAVE_WDATA_WIDTH (PORT_CTRL_MMR_SLAVE_WDATA_WIDTH),
      .PORT_CTRL_MMR_SLAVE_BCOUNT_WIDTH (PORT_CTRL_MMR_SLAVE_BCOUNT_WIDTH),
      .PORT_HPS_EMIF_H2E_WIDTH (PORT_HPS_EMIF_H2E_WIDTH),
      .PORT_HPS_EMIF_E2H_WIDTH (PORT_HPS_EMIF_E2H_WIDTH),
      .PORT_HPS_EMIF_H2E_GP_WIDTH (PORT_HPS_EMIF_H2E_GP_WIDTH),
      .PORT_HPS_EMIF_E2H_GP_WIDTH (PORT_HPS_EMIF_E2H_GP_WIDTH),
      .PORT_CAL_DEBUG_ADDRESS_WIDTH (PORT_CAL_DEBUG_ADDRESS_WIDTH),
      .PORT_CAL_DEBUG_RDATA_WIDTH (PORT_CAL_DEBUG_RDATA_WIDTH),
      .PORT_CAL_DEBUG_WDATA_WIDTH (PORT_CAL_DEBUG_WDATA_WIDTH),
      .PORT_CAL_DEBUG_BYTEEN_WIDTH (PORT_CAL_DEBUG_BYTEEN_WIDTH),
      .PORT_CAL_DEBUG_OUT_ADDRESS_WIDTH (PORT_CAL_DEBUG_OUT_ADDRESS_WIDTH),
      .PORT_CAL_DEBUG_OUT_RDATA_WIDTH (PORT_CAL_DEBUG_OUT_RDATA_WIDTH),
      .PORT_CAL_DEBUG_OUT_WDATA_WIDTH (PORT_CAL_DEBUG_OUT_WDATA_WIDTH),
      .PORT_CAL_DEBUG_OUT_BYTEEN_WIDTH (PORT_CAL_DEBUG_OUT_BYTEEN_WIDTH),
      .PORT_CAL_MASTER_ADDRESS_WIDTH (PORT_CAL_MASTER_ADDRESS_WIDTH),
      .PORT_CAL_MASTER_RDATA_WIDTH (PORT_CAL_MASTER_RDATA_WIDTH),
      .PORT_CAL_MASTER_WDATA_WIDTH (PORT_CAL_MASTER_WDATA_WIDTH),
      .PORT_CAL_MASTER_BYTEEN_WIDTH (PORT_CAL_MASTER_BYTEEN_WIDTH),
      .PORT_DFT_NF_IOAUX_PIO_IN_WIDTH (PORT_DFT_NF_IOAUX_PIO_IN_WIDTH),
      .PORT_DFT_NF_IOAUX_PIO_OUT_WIDTH (PORT_DFT_NF_IOAUX_PIO_OUT_WIDTH),
      .PORT_DFT_NF_PA_DPRIO_REG_ADDR_WIDTH (PORT_DFT_NF_PA_DPRIO_REG_ADDR_WIDTH),
      .PORT_DFT_NF_PA_DPRIO_WRITEDATA_WIDTH (PORT_DFT_NF_PA_DPRIO_WRITEDATA_WIDTH),
      .PORT_DFT_NF_PA_DPRIO_READDATA_WIDTH (PORT_DFT_NF_PA_DPRIO_READDATA_WIDTH),
      .PORT_DFT_NF_PLL_CNTSEL_WIDTH (PORT_DFT_NF_PLL_CNTSEL_WIDTH),
      .PORT_DFT_NF_PLL_NUM_SHIFT_WIDTH (PORT_DFT_NF_PLL_NUM_SHIFT_WIDTH),
      .PORT_DFT_NF_CORE_CLK_BUF_OUT_WIDTH (PORT_DFT_NF_CORE_CLK_BUF_OUT_WIDTH),
      .PORT_DFT_NF_CORE_CLK_LOCKED_WIDTH (PORT_DFT_NF_CORE_CLK_LOCKED_WIDTH),
      .PLL_VCO_FREQ_MHZ_INT (PLL_VCO_FREQ_MHZ_INT),
      .PLL_VCO_TO_MEM_CLK_FREQ_RATIO (PLL_VCO_TO_MEM_CLK_FREQ_RATIO),
      .PLL_PHY_CLK_VCO_PHASE (PLL_PHY_CLK_VCO_PHASE),
      .PLL_VCO_FREQ_PS_STR (PLL_VCO_FREQ_PS_STR),
      .PLL_REF_CLK_FREQ_PS_STR (PLL_REF_CLK_FREQ_PS_STR),
      .PLL_REF_CLK_FREQ_PS (PLL_REF_CLK_FREQ_PS),
      .PLL_SIM_VCO_FREQ_PS (PLL_SIM_VCO_FREQ_PS),
      .PLL_SIM_PHYCLK_0_FREQ_PS (PLL_SIM_PHYCLK_0_FREQ_PS),
      .PLL_SIM_PHYCLK_1_FREQ_PS (PLL_SIM_PHYCLK_1_FREQ_PS),
      .PLL_SIM_PHYCLK_FB_FREQ_PS (PLL_SIM_PHYCLK_FB_FREQ_PS),
      .PLL_SIM_PHY_CLK_VCO_PHASE_PS (PLL_SIM_PHY_CLK_VCO_PHASE_PS),
      .PLL_SIM_CAL_SLAVE_CLK_FREQ_PS (PLL_SIM_CAL_SLAVE_CLK_FREQ_PS),
      .PLL_SIM_CAL_MASTER_CLK_FREQ_PS (PLL_SIM_CAL_MASTER_CLK_FREQ_PS),
      .PLL_M_CNT_HIGH (PLL_M_CNT_HIGH),
      .PLL_M_CNT_LOW (PLL_M_CNT_LOW),
      .PLL_N_CNT_HIGH (PLL_N_CNT_HIGH),
      .PLL_N_CNT_LOW (PLL_N_CNT_LOW),
      .PLL_M_CNT_BYPASS_EN (PLL_M_CNT_BYPASS_EN),
      .PLL_N_CNT_BYPASS_EN (PLL_N_CNT_BYPASS_EN),
      .PLL_M_CNT_EVEN_DUTY_EN (PLL_M_CNT_EVEN_DUTY_EN),
      .PLL_N_CNT_EVEN_DUTY_EN (PLL_N_CNT_EVEN_DUTY_EN),
      .PLL_FBCLK_MUX_1 (PLL_FBCLK_MUX_1),
      .PLL_FBCLK_MUX_2 (PLL_FBCLK_MUX_2),
      .PLL_M_CNT_IN_SRC (PLL_M_CNT_IN_SRC),
      .PLL_CP_SETTING (PLL_CP_SETTING),
      .PLL_BW_CTRL (PLL_BW_CTRL),
      .PLL_BW_SEL (PLL_BW_SEL),
      .PLL_C_CNT_HIGH_0 (PLL_C_CNT_HIGH_0),
      .PLL_C_CNT_LOW_0 (PLL_C_CNT_LOW_0),
      .PLL_C_CNT_PRST_0 (PLL_C_CNT_PRST_0),
      .PLL_C_CNT_PH_MUX_PRST_0 (PLL_C_CNT_PH_MUX_PRST_0),
      .PLL_C_CNT_BYPASS_EN_0 (PLL_C_CNT_BYPASS_EN_0),
      .PLL_C_CNT_EVEN_DUTY_EN_0 (PLL_C_CNT_EVEN_DUTY_EN_0),
      .PLL_C_CNT_FREQ_PS_STR_0 (PLL_C_CNT_FREQ_PS_STR_0),
      .PLL_C_CNT_PHASE_PS_STR_0 (PLL_C_CNT_PHASE_PS_STR_0),
      .PLL_C_CNT_DUTY_CYCLE_0 (PLL_C_CNT_DUTY_CYCLE_0),
      .PLL_C_CNT_OUT_EN_0 (PLL_C_CNT_OUT_EN_0),
      .PLL_C_CNT_HIGH_1 (PLL_C_CNT_HIGH_1),
      .PLL_C_CNT_LOW_1 (PLL_C_CNT_LOW_1),
      .PLL_C_CNT_PRST_1 (PLL_C_CNT_PRST_1),
      .PLL_C_CNT_PH_MUX_PRST_1 (PLL_C_CNT_PH_MUX_PRST_1),
      .PLL_C_CNT_BYPASS_EN_1 (PLL_C_CNT_BYPASS_EN_1),
      .PLL_C_CNT_EVEN_DUTY_EN_1 (PLL_C_CNT_EVEN_DUTY_EN_1),
      .PLL_C_CNT_FREQ_PS_STR_1 (PLL_C_CNT_FREQ_PS_STR_1),
      .PLL_C_CNT_PHASE_PS_STR_1 (PLL_C_CNT_PHASE_PS_STR_1),
      .PLL_C_CNT_DUTY_CYCLE_1 (PLL_C_CNT_DUTY_CYCLE_1),
      .PLL_C_CNT_OUT_EN_1 (PLL_C_CNT_OUT_EN_1),
      .PLL_C_CNT_HIGH_2 (PLL_C_CNT_HIGH_2),
      .PLL_C_CNT_LOW_2 (PLL_C_CNT_LOW_2),
      .PLL_C_CNT_PRST_2 (PLL_C_CNT_PRST_2),
      .PLL_C_CNT_PH_MUX_PRST_2 (PLL_C_CNT_PH_MUX_PRST_2),
      .PLL_C_CNT_BYPASS_EN_2 (PLL_C_CNT_BYPASS_EN_2),
      .PLL_C_CNT_EVEN_DUTY_EN_2 (PLL_C_CNT_EVEN_DUTY_EN_2),
      .PLL_C_CNT_FREQ_PS_STR_2 (PLL_C_CNT_FREQ_PS_STR_2),
      .PLL_C_CNT_PHASE_PS_STR_2 (PLL_C_CNT_PHASE_PS_STR_2),
      .PLL_C_CNT_DUTY_CYCLE_2 (PLL_C_CNT_DUTY_CYCLE_2),
      .PLL_C_CNT_OUT_EN_2 (PLL_C_CNT_OUT_EN_2),
      .PLL_C_CNT_HIGH_3 (PLL_C_CNT_HIGH_3),
      .PLL_C_CNT_LOW_3 (PLL_C_CNT_LOW_3),
      .PLL_C_CNT_PRST_3 (PLL_C_CNT_PRST_3),
      .PLL_C_CNT_PH_MUX_PRST_3 (PLL_C_CNT_PH_MUX_PRST_3),
      .PLL_C_CNT_BYPASS_EN_3 (PLL_C_CNT_BYPASS_EN_3),
      .PLL_C_CNT_EVEN_DUTY_EN_3 (PLL_C_CNT_EVEN_DUTY_EN_3),
      .PLL_C_CNT_FREQ_PS_STR_3 (PLL_C_CNT_FREQ_PS_STR_3),
      .PLL_C_CNT_PHASE_PS_STR_3 (PLL_C_CNT_PHASE_PS_STR_3),
      .PLL_C_CNT_DUTY_CYCLE_3 (PLL_C_CNT_DUTY_CYCLE_3),
      .PLL_C_CNT_OUT_EN_3 (PLL_C_CNT_OUT_EN_3),
      .PLL_C_CNT_HIGH_4 (PLL_C_CNT_HIGH_4),
      .PLL_C_CNT_LOW_4 (PLL_C_CNT_LOW_4),
      .PLL_C_CNT_PRST_4 (PLL_C_CNT_PRST_4),
      .PLL_C_CNT_PH_MUX_PRST_4 (PLL_C_CNT_PH_MUX_PRST_4),
      .PLL_C_CNT_BYPASS_EN_4 (PLL_C_CNT_BYPASS_EN_4),
      .PLL_C_CNT_EVEN_DUTY_EN_4 (PLL_C_CNT_EVEN_DUTY_EN_4),
      .PLL_C_CNT_FREQ_PS_STR_4 (PLL_C_CNT_FREQ_PS_STR_4),
      .PLL_C_CNT_PHASE_PS_STR_4 (PLL_C_CNT_PHASE_PS_STR_4),
      .PLL_C_CNT_DUTY_CYCLE_4 (PLL_C_CNT_DUTY_CYCLE_4),
      .PLL_C_CNT_OUT_EN_4 (PLL_C_CNT_OUT_EN_4),
      .PLL_C_CNT_HIGH_5 (PLL_C_CNT_HIGH_5),
      .PLL_C_CNT_LOW_5 (PLL_C_CNT_LOW_5),
      .PLL_C_CNT_PRST_5 (PLL_C_CNT_PRST_5),
      .PLL_C_CNT_PH_MUX_PRST_5 (PLL_C_CNT_PH_MUX_PRST_5),
      .PLL_C_CNT_BYPASS_EN_5 (PLL_C_CNT_BYPASS_EN_5),
      .PLL_C_CNT_EVEN_DUTY_EN_5 (PLL_C_CNT_EVEN_DUTY_EN_5),
      .PLL_C_CNT_FREQ_PS_STR_5 (PLL_C_CNT_FREQ_PS_STR_5),
      .PLL_C_CNT_PHASE_PS_STR_5 (PLL_C_CNT_PHASE_PS_STR_5),
      .PLL_C_CNT_DUTY_CYCLE_5 (PLL_C_CNT_DUTY_CYCLE_5),
      .PLL_C_CNT_OUT_EN_5 (PLL_C_CNT_OUT_EN_5),
      .PLL_C_CNT_HIGH_6 (PLL_C_CNT_HIGH_6),
      .PLL_C_CNT_LOW_6 (PLL_C_CNT_LOW_6),
      .PLL_C_CNT_PRST_6 (PLL_C_CNT_PRST_6),
      .PLL_C_CNT_PH_MUX_PRST_6 (PLL_C_CNT_PH_MUX_PRST_6),
      .PLL_C_CNT_BYPASS_EN_6 (PLL_C_CNT_BYPASS_EN_6),
      .PLL_C_CNT_EVEN_DUTY_EN_6 (PLL_C_CNT_EVEN_DUTY_EN_6),
      .PLL_C_CNT_FREQ_PS_STR_6 (PLL_C_CNT_FREQ_PS_STR_6),
      .PLL_C_CNT_PHASE_PS_STR_6 (PLL_C_CNT_PHASE_PS_STR_6),
      .PLL_C_CNT_DUTY_CYCLE_6 (PLL_C_CNT_DUTY_CYCLE_6),
      .PLL_C_CNT_OUT_EN_6 (PLL_C_CNT_OUT_EN_6),
      .PLL_C_CNT_HIGH_7 (PLL_C_CNT_HIGH_7),
      .PLL_C_CNT_LOW_7 (PLL_C_CNT_LOW_7),
      .PLL_C_CNT_PRST_7 (PLL_C_CNT_PRST_7),
      .PLL_C_CNT_PH_MUX_PRST_7 (PLL_C_CNT_PH_MUX_PRST_7),
      .PLL_C_CNT_BYPASS_EN_7 (PLL_C_CNT_BYPASS_EN_7),
      .PLL_C_CNT_EVEN_DUTY_EN_7 (PLL_C_CNT_EVEN_DUTY_EN_7),
      .PLL_C_CNT_FREQ_PS_STR_7 (PLL_C_CNT_FREQ_PS_STR_7),
      .PLL_C_CNT_PHASE_PS_STR_7 (PLL_C_CNT_PHASE_PS_STR_7),
      .PLL_C_CNT_DUTY_CYCLE_7 (PLL_C_CNT_DUTY_CYCLE_7),
      .PLL_C_CNT_OUT_EN_7 (PLL_C_CNT_OUT_EN_7),
      .PLL_C_CNT_HIGH_8 (PLL_C_CNT_HIGH_8),
      .PLL_C_CNT_LOW_8 (PLL_C_CNT_LOW_8),
      .PLL_C_CNT_PRST_8 (PLL_C_CNT_PRST_8),
      .PLL_C_CNT_PH_MUX_PRST_8 (PLL_C_CNT_PH_MUX_PRST_8),
      .PLL_C_CNT_BYPASS_EN_8 (PLL_C_CNT_BYPASS_EN_8),
      .PLL_C_CNT_EVEN_DUTY_EN_8 (PLL_C_CNT_EVEN_DUTY_EN_8),
      .PLL_C_CNT_FREQ_PS_STR_8 (PLL_C_CNT_FREQ_PS_STR_8),
      .PLL_C_CNT_PHASE_PS_STR_8 (PLL_C_CNT_PHASE_PS_STR_8),
      .PLL_C_CNT_DUTY_CYCLE_8 (PLL_C_CNT_DUTY_CYCLE_8),
      .PLL_C_CNT_OUT_EN_8 (PLL_C_CNT_OUT_EN_8),
      .SEQ_SYNTH_PARAMS_HEX_FILENAME ("emif_ddr4_ddr4b_altera_emif_arch_nf_170_3eabgiq_seq_params_synth.hex"),
      .SEQ_SIM_PARAMS_HEX_FILENAME ("emif_ddr4_ddr4b_altera_emif_arch_nf_170_3eabgiq_seq_params_sim.hex"),
      .SEQ_CODE_HEX_FILENAME ("emif_ddr4_ddr4b_altera_emif_arch_nf_170_3eabgiq_seq_cal.hex")
   ) arch_inst (
      .global_reset_n (global_reset_n),
      .pll_ref_clk (pll_ref_clk),
      .pll_locked (pll_locked),
      .pll_extra_clk_0 (pll_extra_clk_0),
      .pll_extra_clk_1 (pll_extra_clk_1),
      .pll_extra_clk_2 (pll_extra_clk_2),
      .pll_extra_clk_3 (pll_extra_clk_3),
      .oct_rzqin (oct_rzqin),
      .mem_ck (mem_ck),
      .mem_ck_n (mem_ck_n),
      .mem_a (mem_a),
      .mem_act_n (mem_act_n),
      .mem_ba (mem_ba),
      .mem_bg (mem_bg),
      .mem_c (mem_c),
      .mem_cke (mem_cke),
      .mem_cs_n (mem_cs_n),
      .mem_rm (mem_rm),
      .mem_odt (mem_odt),
      .mem_reset_n (mem_reset_n),
      .mem_par (mem_par),
      .mem_alert_n (mem_alert_n),
      .mem_dqs (mem_dqs),
      .mem_dqs_n (mem_dqs_n),
      .mem_dq (mem_dq),
      .mem_dbi_n (mem_dbi_n),
      .mem_dk (mem_dk),
      .mem_dk_n (mem_dk_n),
      .mem_dka (mem_dka),
      .mem_dka_n (mem_dka_n),
      .mem_dkb (mem_dkb),
      .mem_dkb_n (mem_dkb_n),
      .mem_k (mem_k),
      .mem_k_n (mem_k_n),
      .mem_ras_n (mem_ras_n),
      .mem_cas_n (mem_cas_n),
      .mem_we_n (mem_we_n),
      .mem_ca (mem_ca),
      .mem_ref_n (mem_ref_n),
      .mem_wps_n (mem_wps_n),
      .mem_rps_n (mem_rps_n),
      .mem_doff_n (mem_doff_n),
      .mem_lda_n (mem_lda_n),
      .mem_ldb_n (mem_ldb_n),
      .mem_rwa_n (mem_rwa_n),
      .mem_rwb_n (mem_rwb_n),
      .mem_lbk0_n (mem_lbk0_n),
      .mem_lbk1_n (mem_lbk1_n),
      .mem_cfg_n (mem_cfg_n),
      .mem_ap (mem_ap),
      .mem_ainv (mem_ainv),
      .mem_dm (mem_dm),
      .mem_bws_n (mem_bws_n),
      .mem_d (mem_d),
      .mem_dqa (mem_dqa),
      .mem_dqb (mem_dqb),
      .mem_dinva (mem_dinva),
      .mem_dinvb (mem_dinvb),
      .mem_q (mem_q),
      .mem_qk (mem_qk),
      .mem_qk_n (mem_qk_n),
      .mem_qka (mem_qka),
      .mem_qka_n (mem_qka_n),
      .mem_qkb (mem_qkb),
      .mem_qkb_n (mem_qkb_n),
      .mem_cq (mem_cq),
      .mem_cq_n (mem_cq_n),
      .mem_pe_n (mem_pe_n),
      .local_cal_success (local_cal_success),
      .local_cal_fail (local_cal_fail),
      .vid_cal_done_persist (vid_cal_done_persist),
      .afi_reset_n (afi_reset_n),
      .afi_clk (afi_clk),
      .afi_half_clk (afi_half_clk),
      .emif_usr_reset_n (emif_usr_reset_n),
      .emif_usr_clk (emif_usr_clk),
      .emif_usr_half_clk (emif_usr_half_clk),
      .emif_usr_reset_n_sec (emif_usr_reset_n_sec),
      .emif_usr_clk_sec (emif_usr_clk_sec),
      .emif_usr_half_clk_sec (emif_usr_half_clk_sec),
      .cal_master_reset_n (cal_master_reset_n),
      .cal_master_clk (cal_master_clk),
      .cal_slave_reset_n (cal_slave_reset_n),
      .cal_slave_clk (cal_slave_clk),
      .cal_slave_reset_n_in (cal_slave_reset_n_in),
      .cal_slave_clk_in (cal_slave_clk_in),
      .cal_debug_reset_n (cal_debug_reset_n),
      .cal_debug_clk (cal_debug_clk),
      .cal_debug_out_reset_n (cal_debug_out_reset_n),
      .cal_debug_out_clk (cal_debug_out_clk),
      .clks_sharing_master_out (clks_sharing_master_out),
      .clks_sharing_slave_in (clks_sharing_slave_in),
      .afi_cal_success (afi_cal_success),
      .afi_cal_fail (afi_cal_fail),
      .afi_cal_req (afi_cal_req),
      .afi_rlat (afi_rlat),
      .afi_wlat (afi_wlat),
      .afi_seq_busy (afi_seq_busy),
      .afi_ctl_refresh_done (afi_ctl_refresh_done),
      .afi_ctl_long_idle (afi_ctl_long_idle),
      .afi_mps_req (afi_mps_req),
      .afi_mps_ack (afi_mps_ack),
      .afi_addr (afi_addr),
      .afi_ba (afi_ba),
      .afi_bg (afi_bg),
      .afi_c (afi_c),
      .afi_cke (afi_cke),
      .afi_cs_n (afi_cs_n),
      .afi_rm (afi_rm),
      .afi_odt (afi_odt),
      .afi_ras_n (afi_ras_n),
      .afi_cas_n (afi_cas_n),
      .afi_we_n (afi_we_n),
      .afi_rst_n (afi_rst_n),
      .afi_act_n (afi_act_n),
      .afi_par (afi_par),
      .afi_ca (afi_ca),
      .afi_ref_n (afi_ref_n),
      .afi_wps_n (afi_wps_n),
      .afi_rps_n (afi_rps_n),
      .afi_doff_n (afi_doff_n),
      .afi_ld_n (afi_ld_n),
      .afi_rw_n (afi_rw_n),
      .afi_lbk0_n (afi_lbk0_n),
      .afi_lbk1_n (afi_lbk1_n),
      .afi_cfg_n (afi_cfg_n),
      .afi_ap (afi_ap),
      .afi_ainv (afi_ainv),
      .afi_dm (afi_dm),
      .afi_dm_n (afi_dm_n),
      .afi_bws_n (afi_bws_n),
      .afi_rdata_dbi_n (afi_rdata_dbi_n),
      .afi_wdata_dbi_n (afi_wdata_dbi_n),
      .afi_rdata_dinv (afi_rdata_dinv),
      .afi_wdata_dinv (afi_wdata_dinv),
      .afi_dqs_burst (afi_dqs_burst),
      .afi_wdata_valid (afi_wdata_valid),
      .afi_wdata (afi_wdata),
      .afi_rdata_en_full (afi_rdata_en_full),
      .afi_rdata (afi_rdata),
      .afi_rdata_valid (afi_rdata_valid),
      .afi_rrank (afi_rrank),
      .afi_wrank (afi_wrank),
      .afi_alert_n (afi_alert_n),
      .afi_pe_n (afi_pe_n),
      .ast_cmd_data_0 (ast_cmd_data_0),
      .ast_cmd_valid_0 (ast_cmd_valid_0),
      .ast_cmd_ready_0 (ast_cmd_ready_0),
      .ast_cmd_data_1 (ast_cmd_data_1),
      .ast_cmd_valid_1 (ast_cmd_valid_1),
      .ast_cmd_ready_1 (ast_cmd_ready_1),
      .ast_wr_data_0 (ast_wr_data_0),
      .ast_wr_valid_0 (ast_wr_valid_0),
      .ast_wr_ready_0 (ast_wr_ready_0),
      .ast_wr_data_1 (ast_wr_data_1),
      .ast_wr_valid_1 (ast_wr_valid_1),
      .ast_wr_ready_1 (ast_wr_ready_1),
      .ast_rd_data_0 (ast_rd_data_0),
      .ast_rd_valid_0 (ast_rd_valid_0),
      .ast_rd_ready_0 (ast_rd_ready_0),
      .ast_rd_data_1 (ast_rd_data_1),
      .ast_rd_valid_1 (ast_rd_valid_1),
      .ast_rd_ready_1 (ast_rd_ready_1),
      .amm_ready_0 (amm_ready_0),
      .amm_read_0 (amm_read_0),
      .amm_write_0 (amm_write_0),
      .amm_address_0 (amm_address_0),
      .amm_readdata_0 (amm_readdata_0),
      .amm_writedata_0 (amm_writedata_0),
      .amm_burstcount_0 (amm_burstcount_0),
      .amm_byteenable_0 (amm_byteenable_0),
      .amm_beginbursttransfer_0 (amm_beginbursttransfer_0),
      .amm_readdatavalid_0 (amm_readdatavalid_0),
      .amm_ready_1 (amm_ready_1),
      .amm_read_1 (amm_read_1),
      .amm_write_1 (amm_write_1),
      .amm_address_1 (amm_address_1),
      .amm_readdata_1 (amm_readdata_1),
      .amm_writedata_1 (amm_writedata_1),
      .amm_burstcount_1 (amm_burstcount_1),
      .amm_byteenable_1 (amm_byteenable_1),
      .amm_beginbursttransfer_1 (amm_beginbursttransfer_1),
      .amm_readdatavalid_1 (amm_readdatavalid_1),
      .ctrl_user_priority_hi_0 (ctrl_user_priority_hi_0),
      .ctrl_user_priority_hi_1 (ctrl_user_priority_hi_1),
      .ctrl_auto_precharge_req_0 (ctrl_auto_precharge_req_0),
      .ctrl_auto_precharge_req_1 (ctrl_auto_precharge_req_1),
      .ctrl_user_refresh_req (ctrl_user_refresh_req),
      .ctrl_user_refresh_bank (ctrl_user_refresh_bank),
      .ctrl_user_refresh_ack (ctrl_user_refresh_ack),
      .ctrl_self_refresh_req (ctrl_self_refresh_req),
      .ctrl_self_refresh_ack (ctrl_self_refresh_ack),
      .ctrl_will_refresh (ctrl_will_refresh),
      .ctrl_deep_power_down_req (ctrl_deep_power_down_req),
      .ctrl_deep_power_down_ack (ctrl_deep_power_down_ack),
      .ctrl_power_down_ack (ctrl_power_down_ack),
      .ctrl_zq_cal_long_req (ctrl_zq_cal_long_req),
      .ctrl_zq_cal_short_req (ctrl_zq_cal_short_req),
      .ctrl_zq_cal_ack (ctrl_zq_cal_ack),
      .ctrl_ecc_write_info_0 (ctrl_ecc_write_info_0),
      .ctrl_ecc_rdata_id_0 (ctrl_ecc_rdata_id_0),
      .ctrl_ecc_read_info_0 (ctrl_ecc_read_info_0),
      .ctrl_ecc_cmd_info_0 (ctrl_ecc_cmd_info_0),
      .ctrl_ecc_idle_0 (ctrl_ecc_idle_0),
      .ctrl_ecc_wr_pointer_info_0 (ctrl_ecc_wr_pointer_info_0),
      .ctrl_ecc_write_info_1 (ctrl_ecc_write_info_1),
      .ctrl_ecc_rdata_id_1 (ctrl_ecc_rdata_id_1),
      .ctrl_ecc_read_info_1 (ctrl_ecc_read_info_1),
      .ctrl_ecc_cmd_info_1 (ctrl_ecc_cmd_info_1),
      .ctrl_ecc_idle_1 (ctrl_ecc_idle_1),
      .ctrl_ecc_wr_pointer_info_1 (ctrl_ecc_wr_pointer_info_1),
      .mmr_slave_waitrequest_0 (mmr_slave_waitrequest_0),
      .mmr_slave_read_0 (mmr_slave_read_0),
      .mmr_slave_write_0 (mmr_slave_write_0),
      .mmr_slave_address_0 (mmr_slave_address_0),
      .mmr_slave_readdata_0 (mmr_slave_readdata_0),
      .mmr_slave_writedata_0 (mmr_slave_writedata_0),
      .mmr_slave_burstcount_0 (mmr_slave_burstcount_0),
      .mmr_slave_beginbursttransfer_0 (mmr_slave_beginbursttransfer_0),
      .mmr_slave_readdatavalid_0 (mmr_slave_readdatavalid_0),
      .mmr_slave_waitrequest_1 (mmr_slave_waitrequest_1),
      .mmr_slave_read_1 (mmr_slave_read_1),
      .mmr_slave_write_1 (mmr_slave_write_1),
      .mmr_slave_address_1 (mmr_slave_address_1),
      .mmr_slave_readdata_1 (mmr_slave_readdata_1),
      .mmr_slave_writedata_1 (mmr_slave_writedata_1),
      .mmr_slave_burstcount_1 (mmr_slave_burstcount_1),
      .mmr_slave_beginbursttransfer_1 (mmr_slave_beginbursttransfer_1),
      .mmr_slave_readdatavalid_1 (mmr_slave_readdatavalid_1),
      .hps_to_emif (hps_to_emif),
      .emif_to_hps (emif_to_hps),
      .hps_to_emif_gp (hps_to_emif_gp),
      .emif_to_hps_gp (emif_to_hps_gp),
      .cal_debug_waitrequest (cal_debug_waitrequest),
      .cal_debug_read (cal_debug_read),
      .cal_debug_write (cal_debug_write),
      .cal_debug_addr (cal_debug_addr),
      .cal_debug_read_data (cal_debug_read_data),
      .cal_debug_write_data (cal_debug_write_data),
      .cal_debug_byteenable (cal_debug_byteenable),
      .cal_debug_read_data_valid (cal_debug_read_data_valid),
      .cal_debug_out_waitrequest (cal_debug_out_waitrequest),
      .cal_debug_out_read (cal_debug_out_read),
      .cal_debug_out_write (cal_debug_out_write),
      .cal_debug_out_addr (cal_debug_out_addr),
      .cal_debug_out_read_data (cal_debug_out_read_data),
      .cal_debug_out_write_data (cal_debug_out_write_data),
      .cal_debug_out_byteenable (cal_debug_out_byteenable),
      .cal_debug_out_read_data_valid (cal_debug_out_read_data_valid),
      .cal_master_waitrequest (cal_master_waitrequest),
      .cal_master_read (cal_master_read),
      .cal_master_write (cal_master_write),
      .cal_master_addr (cal_master_addr),
      .cal_master_read_data (cal_master_read_data),
      .cal_master_write_data (cal_master_write_data),
      .cal_master_byteenable (cal_master_byteenable),
      .cal_master_read_data_valid (cal_master_read_data_valid),
      .cal_master_burstcount (cal_master_burstcount),
      .cal_master_debugaccess (cal_master_debugaccess),
      .ioaux_pio_in (ioaux_pio_in),
      .ioaux_pio_out (ioaux_pio_out),
      .pa_dprio_clk (pa_dprio_clk),
      .pa_dprio_read (pa_dprio_read),
      .pa_dprio_reg_addr (pa_dprio_reg_addr),
      .pa_dprio_rst_n (pa_dprio_rst_n),
      .pa_dprio_write (pa_dprio_write),
      .pa_dprio_writedata (pa_dprio_writedata),
      .pa_dprio_block_select (pa_dprio_block_select),
      .pa_dprio_readdata (pa_dprio_readdata),
      .pll_phase_en (pll_phase_en),
      .pll_up_dn (pll_up_dn),
      .pll_cnt_sel (pll_cnt_sel),
      .pll_num_phase_shifts (pll_num_phase_shifts),
      .pll_phase_done (pll_phase_done),
      .dft_core_clk_buf_out (dft_core_clk_buf_out),
      .dft_core_clk_locked (dft_core_clk_locked)
   );
endmodule
