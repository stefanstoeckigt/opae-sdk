// ddr4b_clock_bridge.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module ddr4b_clock_bridge (
		input  wire  in_clk,  //  in_clk.clk
		output wire  out_clk  // out_clk.clk
	);

	assign out_clk = in_clk;

endmodule
